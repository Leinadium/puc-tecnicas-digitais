CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 200 5 150 10
2 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
170 176 283 273
42991634 0
0
6 Title:
5 Name:
0
0
0
169
9 Terminal~
194 166 486 0 1 3
0 5
0
0 0 49504 270
6 nclock
2 -4 44 4
3 T83
-10 -32 11 -24
0
7 nclock;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3901 0 0
2
44519.5 0
0
13 Logic Switch~
5 1668 296 0 1 11
0 51
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6295 0 0
2
5.90009e-315 0
0
13 Logic Switch~
5 2475 189 0 1 11
0 64
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
332 0 0
2
5.90009e-315 5.43969e-315
0
13 Logic Switch~
5 2470 331 0 1 11
0 62
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9737 0 0
2
5.90009e-315 5.4371e-315
0
13 Logic Switch~
5 2472 479 0 1 11
0 60
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9910 0 0
2
5.90009e-315 5.43451e-315
0
13 Logic Switch~
5 2475 619 0 1 11
0 58
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3834 0 0
2
5.90009e-315 5.43192e-315
0
13 Logic Switch~
5 2410 149 0 1 11
0 56
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3138 0 0
2
5.90009e-315 5.42933e-315
0
13 Logic Switch~
5 1596 154 0 10 11
0 52 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5409 0 0
2
5.90009e-315 0
0
9 Inverter~
13 1326 1504 0 2 22
0 3 41
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
983 0 0
2
44519.5 0
0
9 Terminal~
194 1438 1486 0 1 3
0 2
0
0 0 49520 0
4 orup
-14 -22 14 -14
3 T82
-11 -32 10 -24
0
5 orup;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
6652 0 0
2
44519.5 3
0
9 Terminal~
194 1267 1493 0 1 3
0 3
0
0 0 49520 0
7 qquatro
-24 -22 25 -14
3 T81
-11 -32 10 -24
0
8 qquatro;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
4281 0 0
2
44519.5 2
0
9 Terminal~
194 1304 1477 0 1 3
0 4
0
0 0 49520 0
6 clockd
-20 -22 22 -14
3 T80
-11 -32 10 -24
0
7 clockd;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
6847 0 0
2
44519.5 1
0
5 4081~
219 1386 1495 0 3 22
0 4 41 2
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U16B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 7 0
1 U
6543 0 0
2
44519.5 0
0
5 4081~
219 1082 1495 0 3 22
0 5 3 2
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U16A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 7 0
1 U
7168 0 0
2
44519.5 3
0
9 Terminal~
194 1000 1477 0 1 3
0 5
0
0 0 49520 0
5 clock
-17 -22 18 -14
3 T77
-11 -32 10 -24
0
6 clock;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
3828 0 0
2
44519.5 2
0
9 Terminal~
194 1035 1494 0 1 3
0 3
0
0 0 49520 0
7 qquatro
-24 -22 25 -14
3 T78
-11 -32 10 -24
0
8 qquatro;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
955 0 0
2
44519.5 1
0
9 Terminal~
194 1134 1486 0 1 3
0 2
0
0 0 49520 0
4 orup
-14 -22 14 -14
3 T79
-11 -32 10 -24
0
5 orup;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
7782 0 0
2
44519.5 0
0
5 4013~
219 1710 1295 0 6 22
0 9 42 6 7 78 8
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U18B
21 -54 49 -46
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 9 0
1 U
824 0 0
2
44519.5 5
0
2 +V
167 1649 1247 0 1 3
0 42
0
0 0 54256 0
3 10V
-11 -22 10 -14
3 V18
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6983 0 0
2
44519.5 4
0
9 Terminal~
194 1609 1266 0 1 3
0 6
0
0 0 49520 0
4 ddup
-14 -22 14 -14
3 T72
-11 -32 10 -24
0
5 ddup;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
3185 0 0
2
44519.5 3
0
9 Terminal~
194 1642 1304 0 1 3
0 7
0
0 0 49520 0
6 dddown
-21 -21 21 -13
3 T71
-11 -32 10 -24
0
7 dddown;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
4213 0 0
2
44519.5 2
0
9 Terminal~
194 1792 1249 0 1 3
0 8
0
0 0 49520 0
5 ddout
-17 -22 18 -14
3 T70
-11 -32 10 -24
0
6 ddout;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
9765 0 0
2
44519.5 1
0
7 Ground~
168 1681 1337 0 1 3
0 9
0
0 0 53360 0
0
5 GND22
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8986 0 0
2
44519.5 0
0
5 4013~
219 1400 1295 0 6 22
0 9 43 2 10 79 11
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U18A
21 -54 49 -46
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 9 0
1 U
3273 0 0
2
44519.5 5
0
2 +V
167 1339 1247 0 1 3
0 43
0
0 0 54256 0
3 10V
-11 -22 10 -14
3 V17
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5636 0 0
2
44519.5 4
0
9 Terminal~
194 1299 1266 0 1 3
0 2
0
0 0 49520 0
4 orup
-14 -22 14 -14
3 T69
-11 -32 10 -24
0
5 orup;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
327 0 0
2
44519.5 3
0
9 Terminal~
194 1332 1304 0 1 3
0 10
0
0 0 49520 0
6 ordown
-21 -22 21 -14
3 T68
-11 -32 10 -24
0
7 ordown;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
9233 0 0
2
44519.5 2
0
9 Terminal~
194 1482 1249 0 1 3
0 11
0
0 0 49520 0
5 orout
-17 -22 18 -14
3 T67
-11 -32 10 -24
0
6 orout;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
3875 0 0
2
44519.5 1
0
7 Ground~
168 1371 1337 0 1 3
0 9
0
0 0 53360 0
0
5 GND21
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9991 0 0
2
44519.5 0
0
9 Terminal~
194 1792 1033 0 1 3
0 3
0
0 0 49520 0
7 qquatro
-24 -22 25 -14
3 T76
-11 -32 10 -24
0
8 qquatro;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
3221 0 0
2
44519.5 0
0
7 Ground~
168 1076 1338 0 1 3
0 9
0
0 0 53360 0
0
5 GND23
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8874 0 0
2
44519.5 0
0
9 Terminal~
194 1187 1250 0 1 3
0 12
0
0 0 49520 0
4 wout
-14 -22 14 -14
3 T75
-11 -32 10 -24
0
5 wout;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
7400 0 0
2
44519.5 0
0
9 Terminal~
194 1037 1305 0 1 3
0 13
0
0 0 49520 0
5 wdown
-18 -22 17 -14
3 T74
-11 -32 10 -24
0
6 wdown;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
3623 0 0
2
44519.5 0
0
9 Terminal~
194 1004 1267 0 1 3
0 14
0
0 0 49520 0
3 wup
-11 -22 10 -14
3 T73
-11 -32 10 -24
0
4 wup;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
3311 0 0
2
44519.5 0
0
2 +V
167 1044 1248 0 1 3
0 44
0
0 0 54256 0
3 10V
-11 -22 10 -14
3 V16
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5736 0 0
2
44519.5 0
0
5 4013~
219 1105 1296 0 6 22
0 9 44 14 13 80 12
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U17B
21 -54 49 -46
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 8 0
1 U
3143 0 0
2
44519.5 0
0
7 Ground~
168 1645 1117 0 1 3
0 9
0
0 0 53360 0
0
5 GND20
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5835 0 0
2
44519.4 4
0
2 +V
167 1620 942 0 1 3
0 45
0
0 0 54256 0
3 10V
-11 -22 10 -14
3 V11
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5108 0 0
2
44519.4 3
0
9 Terminal~
194 1600 994 0 1 3
0 15
0
0 0 49520 0
6 pqdown
-22 -22 20 -14
3 T66
-11 -32 10 -24
0
7 pqdown;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
3320 0 0
2
44519.4 2
0
9 Terminal~
194 1639 988 0 1 3
0 16
0
0 0 49520 0
4 pqup
-15 -22 13 -14
3 T65
-11 -32 10 -24
0
5 pqup;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
523 0 0
2
44519.4 1
0
7 74LS193
137 1693 1024 0 14 29
0 16 15 45 9 9 9 9 9 81
82 83 3 84 85
0
0 0 4848 0
7 74LS193
-24 -51 25 -43
3 U15
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 0 0 0 0
1 U
3557 0 0
2
44519.4 0
0
7 74LS193
137 1374 1025 0 14 29
0 17 9 46 9 9 9 9 9 86
87 88 89 90 91
0
0 0 4848 0
7 74LS193
-24 -51 25 -43
3 U14
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 0 0 0 0
1 U
7246 0 0
2
44519.4 3
0
7 Ground~
168 1325 1113 0 1 3
0 9
0
0 0 53360 0
0
5 GND19
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3916 0 0
2
44519.4 2
0
2 +V
167 1292 955 0 1 3
0 46
0
0 0 54256 0
3 10V
-11 -22 10 -14
3 V10
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
614 0 0
2
44519.4 1
0
9 Terminal~
194 1260 989 0 1 3
0 17
0
0 0 49520 0
7 pinicio
-25 -22 24 -14
3 T63
-11 -32 10 -24
0
8 pinicio;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
8494 0 0
2
44519.4 0
0
7 Ground~
168 1904 302 0 1 3
0 9
0
0 0 53360 0
0
5 GND18
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
774 0 0
2
5.90009e-315 0
0
5 4013~
219 2541 225 0 6 22
0 9 64 56 9 92 63
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U10A
23 -61 51 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 5 0
1 U
715 0 0
2
5.90009e-315 5.42414e-315
0
7 Ground~
168 2647 149 0 1 3
0 9
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3281 0 0
2
5.90009e-315 5.41896e-315
0
7 Ground~
168 2541 249 0 1 3
0 9
0
0 0 53360 0
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3593 0 0
2
5.90009e-315 5.41378e-315
0
14 Logic Display~
6 2611 171 0 1 2
10 63
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7233 0 0
2
5.90009e-315 5.4086e-315
0
14 Logic Display~
6 2610 313 0 1 2
10 61
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3410 0 0
2
5.90009e-315 5.40342e-315
0
7 Ground~
168 2538 393 0 1 3
0 9
0
0 0 53360 0
0
5 GND11
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3616 0 0
2
5.90009e-315 5.39824e-315
0
7 Ground~
168 2645 290 0 1 3
0 9
0
0 0 53360 0
0
5 GND12
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5202 0 0
2
5.90009e-315 5.39306e-315
0
5 4013~
219 2538 367 0 6 22
0 9 62 56 9 93 61
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U10B
23 -61 51 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 5 0
1 U
9145 0 0
2
5.90009e-315 5.38788e-315
0
14 Logic Display~
6 2608 461 0 1 2
10 59
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9815 0 0
2
5.90009e-315 5.37752e-315
0
7 Ground~
168 2538 539 0 1 3
0 9
0
0 0 53360 0
0
5 GND13
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4766 0 0
2
5.90009e-315 5.36716e-315
0
7 Ground~
168 2645 434 0 1 3
0 9
0
0 0 53360 0
0
5 GND14
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8325 0 0
2
5.90009e-315 5.3568e-315
0
5 4013~
219 2538 515 0 6 22
0 9 60 56 9 94 59
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U11A
23 -61 51 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 6 0
1 U
7196 0 0
2
5.90009e-315 5.34643e-315
0
14 Logic Display~
6 2611 601 0 1 2
10 57
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3567 0 0
2
5.90009e-315 5.32571e-315
0
7 Ground~
168 2541 679 0 1 3
0 9
0
0 0 53360 0
0
5 GND15
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5877 0 0
2
5.90009e-315 5.30499e-315
0
7 Ground~
168 2641 578 0 1 3
0 9
0
0 0 53360 0
0
5 GND16
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4785 0 0
2
5.90009e-315 5.26354e-315
0
5 4013~
219 2541 655 0 6 22
0 9 58 56 9 95 57
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U11B
23 -61 51 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 6 0
1 U
3822 0 0
2
5.90009e-315 0
0
7 74LS245
64 1959 312 0 18 37
0 96 97 98 99 53 54 55 65 100
101 102 103 47 48 49 50 9 52
0
0 0 4848 0
7 74LS245
-24 -60 25 -52
3 U13
-11 -61 10 -53
0
16 DVCC=20;DGND=10;
192 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i]
+ [%20bi %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP14
37

0 9 8 7 6 5 4 3 2 11
12 13 14 15 16 17 18 19 1 9
8 7 6 5 4 3 2 11 12 13
14 15 16 17 18 19 1 0
65 0 0 512 1 0 0 0
1 U
7640 0 0
2
5.90009e-315 0
0
7 Ground~
168 1624 479 0 1 3
0 9
0
0 0 53360 0
0
5 GND17
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9221 0 0
2
5.90009e-315 0
0
6 1K RAM
79 1672 404 0 20 41
0 9 9 9 9 9 9 66 67 68
69 104 105 106 107 53 54 55 65 51
52
0
0 0 4848 0
5 RAM1K
-17 -19 18 -11
3 U12
-11 -70 10 -62
0
16 DVCC=22;DGND=11;
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 512 1 0 0 0
1 U
6484 0 0
2
5.90009e-315 0
0
8 Hex Key~
166 1246 304 0 11 12
0 69 68 67 66 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3689 0 0
2
5.90009e-315 0
0
9 Inverter~
13 762 176 0 2 22
0 32 70
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
3952 0 0
2
44519.4 0
0
9 Terminal~
194 775 217 0 1 3
0 5
0
0 0 49520 180
5 clock
6 -7 41 1
3 T64
-10 -32 11 -24
0
6 clock;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3631 0 0
2
44519.4 1
0
9 2-In AND~
219 821 185 0 3 22
0 70 5 33
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
9359 0 0
2
44519.4 2
0
9 Terminal~
194 86 218 0 1 3
0 18
0
0 0 49520 180
7 output3
-46 4 3 12
3 T60
-10 -32 11 -24
0
8 output3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5584 0 0
2
44519.4 3
0
12 Hex Display~
7 89 179 0 16 19
10 19 20 18 21 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4973 0 0
2
44519.4 4
0
9 Terminal~
194 98 218 0 1 3
0 19
0
0 0 49520 180
7 output1
7 -11 56 -3
3 T57
-10 -32 11 -24
0
8 output1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3239 0 0
2
44519.4 5
0
9 Terminal~
194 92 218 0 1 3
0 20
0
0 0 49520 180
7 output2
3 5 52 13
3 T58
-10 -32 11 -24
0
8 output2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4244 0 0
2
44519.4 6
0
9 Terminal~
194 80 218 0 1 3
0 21
0
0 0 49520 180
7 output4
-56 -9 -7 -1
3 T59
-10 -32 11 -24
0
8 output4;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3391 0 0
2
44519.4 7
0
6 74LS83
105 547 569 0 14 29
0 9 9 30 25 9 22 71 24 9
26 27 29 28 108
0
0 0 4848 0
6 74LS83
-21 -60 21 -52
2 U4
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
4243 0 0
2
44519.4 8
0
9 Inverter~
13 420 587 0 2 22
0 23 71
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3907 0 0
2
44519.4 9
0
9 Terminal~
194 489 580 0 1 3
0 22
0
0 0 49520 90
6 linha1
-52 -7 -10 1
3 T23
-10 -32 11 -24
0
7 linha1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
728 0 0
2
44519.4 10
0
9 Terminal~
194 393 589 0 1 3
0 23
0
0 0 49520 90
6 linha3
-52 -7 -10 1
3 T24
-10 -32 11 -24
0
7 linha3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3585 0 0
2
44519.4 11
0
9 Terminal~
194 489 598 0 1 3
0 24
0
0 0 49520 90
6 linha2
-52 -7 -10 1
3 T25
-10 -32 11 -24
0
7 linha2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3565 0 0
2
44519.4 12
0
7 Ground~
168 506 635 0 1 3
0 9
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3966 0 0
2
44519.4 13
0
9 Terminal~
194 483 562 0 1 3
0 25
0
0 0 49520 90
6 clock2
-48 -6 -6 2
3 T26
-10 -32 11 -24
0
7 clock2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3714 0 0
2
44519.4 14
0
9 Terminal~
194 616 561 0 1 3
0 26
0
0 0 49520 270
3 sn3
12 -4 33 4
3 T30
-10 -32 11 -24
0
4 sn3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3406 0 0
2
44519.4 15
0
9 Terminal~
194 616 570 0 1 3
0 27
0
0 0 49520 270
3 sn2
12 -4 33 4
3 T31
-10 -32 11 -24
0
4 sn2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3132 0 0
2
44519.4 16
0
9 Terminal~
194 616 588 0 1 3
0 28
0
0 0 49520 270
3 sn0
12 -4 33 4
3 T32
-10 -32 11 -24
0
4 sn0;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3842 0 0
2
44519.4 17
0
9 Terminal~
194 616 579 0 1 3
0 29
0
0 0 49520 270
3 sn1
12 -4 33 4
3 T33
-10 -32 11 -24
0
4 sn1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6183 0 0
2
44519.4 18
0
9 Terminal~
194 483 553 0 1 3
0 30
0
0 0 49520 90
6 clock3
-48 -6 -6 2
3 T27
-10 -32 11 -24
0
7 clock3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3356 0 0
2
44519.4 19
0
9 Terminal~
194 483 723 0 1 3
0 25
0
0 0 49520 90
6 clock2
-48 -6 -6 2
3 T38
-10 -32 11 -24
0
7 clock2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3525 0 0
2
44519.4 20
0
9 Inverter~
13 516 721 0 2 22
0 25 31
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
3800 0 0
2
44519.4 21
0
9 Terminal~
194 584 713 0 1 3
0 31
0
0 0 49520 270
3 se3
12 -4 33 4
3 T37
-10 -32 11 -24
0
4 se3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
346 0 0
2
44519.4 22
0
9 Terminal~
194 584 722 0 1 3
0 31
0
0 0 49520 270
3 se2
12 -4 33 4
3 T36
-10 -32 11 -24
0
4 se2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3169 0 0
2
44519.4 23
0
9 Terminal~
194 584 740 0 1 3
0 30
0
0 0 49520 270
3 se0
12 -4 33 4
3 T35
-10 -32 11 -24
0
4 se0;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4826 0 0
2
44519.4 24
0
9 Terminal~
194 584 731 0 1 3
0 31
0
0 0 49520 270
3 se1
12 -4 33 4
3 T34
-10 -32 11 -24
0
4 se1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3971 0 0
2
44519.4 25
0
9 Terminal~
194 535 741 0 1 3
0 30
0
0 0 49520 90
6 clock3
-48 -6 -6 2
3 T29
-10 -32 11 -24
0
7 clock3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3607 0 0
2
44519.4 26
0
9 Terminal~
194 166 466 0 1 3
0 5
0
0 0 49520 270
5 clock
5 -4 40 4
3 T28
-10 -32 11 -24
0
6 clock;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3506 0 0
2
44519.4 27
0
9 2-In AND~
219 105 549 0 3 22
0 5 32 72
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
7829 0 0
2
44519.4 28
0
9 Terminal~
194 58 560 0 1 3
0 32
0
0 0 49520 90
5 block
-18 -15 17 -7
3 T62
-10 -32 11 -24
0
6 block;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3890 0 0
2
44519.4 29
0
9 Terminal~
194 777 136 0 1 3
0 32
0
0 0 49520 270
5 block
13 -4 48 4
3 T61
-10 -32 11 -24
0
6 block;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3126 0 0
2
44519.4 30
0
5 4013~
219 974 747 0 6 22
0 9 73 33 9 109 19
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U8B
24 -54 45 -46
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 3 0
1 U
3935 0 0
2
44519.4 31
0
7 Ground~
168 1026 760 0 1 3
0 9
0
0 0 53360 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9746 0 0
2
44519.4 32
0
9 Terminal~
194 1067 712 0 1 3
0 19
0
0 0 49520 270
7 output1
3 -7 52 1
3 T56
-10 -32 11 -24
0
8 output1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7330 0 0
2
44519.4 33
0
9 Terminal~
194 938 731 0 1 3
0 33
0
0 0 49520 90
3 set
-35 -6 -14 2
3 T55
-10 -32 11 -24
0
4 set;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3972 0 0
2
44519.4 34
0
5 4013~
219 971 630 0 6 22
0 9 74 33 9 110 20
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U8A
24 -54 45 -46
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 3 0
1 U
7818 0 0
2
44519.4 35
0
7 Ground~
168 1023 643 0 1 3
0 9
0
0 0 53360 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3818 0 0
2
44519.4 36
0
9 Terminal~
194 1064 595 0 1 3
0 20
0
0 0 49520 270
7 output2
3 -7 52 1
3 T54
-10 -32 11 -24
0
8 output2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8835 0 0
2
44519.4 37
0
9 Terminal~
194 921 614 0 1 3
0 33
0
0 0 49520 90
3 set
-35 -6 -14 2
3 T53
-10 -32 11 -24
0
4 set;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7484 0 0
2
44519.4 38
0
5 4013~
219 968 519 0 6 22
0 9 75 33 9 111 18
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U7B
24 -54 45 -46
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 2 0
1 U
792 0 0
2
44519.4 39
0
7 Ground~
168 1020 532 0 1 3
0 9
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3826 0 0
2
44519.4 40
0
9 Terminal~
194 1061 484 0 1 3
0 18
0
0 0 49520 270
7 output3
3 -7 52 1
3 T52
-10 -32 11 -24
0
8 output3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7958 0 0
2
44519.4 41
0
9 Terminal~
194 920 503 0 1 3
0 33
0
0 0 49520 90
3 set
-35 -6 -14 2
3 T49
-10 -32 11 -24
0
4 set;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6736 0 0
2
44519.4 42
0
9 Terminal~
194 912 390 0 1 3
0 33
0
0 0 49520 90
3 set
-35 -6 -14 2
3 T51
-10 -32 11 -24
0
4 set;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3755 0 0
2
44519.4 43
0
9 Terminal~
194 872 186 0 1 3
0 33
0
0 0 49520 270
3 set
12 -4 33 4
3 T50
-10 -32 11 -24
0
4 set;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
397 0 0
2
44519.4 44
0
9 Terminal~
194 1059 371 0 1 3
0 21
0
0 0 49520 270
7 output4
3 -7 52 1
3 T48
-10 -32 11 -24
0
8 output4;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5190 0 0
2
44519.4 45
0
7 Ground~
168 1018 419 0 1 3
0 9
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9188 0 0
2
44519.4 46
0
5 4013~
219 966 406 0 6 22
0 9 76 33 9 112 21
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U7A
24 -54 45 -46
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 2 0
1 U
3651 0 0
2
44519.4 47
0
9 Terminal~
194 741 544 0 1 3
0 34
0
0 0 49520 90
6 linha4
-47 -15 -5 -7
3 T47
-10 -32 11 -24
0
7 linha4;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3415 0 0
2
44519.4 48
0
9 Terminal~
194 741 616 0 1 3
0 30
0
0 0 49520 90
3 se0
-34 -6 -13 2
3 T46
-10 -32 11 -24
0
4 se0;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7597 0 0
2
44519.4 49
0
9 Terminal~
194 741 607 0 1 3
0 28
0
0 0 49520 90
3 sn0
-34 -6 -13 2
3 T45
-10 -32 11 -24
0
4 sn0;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
350 0 0
2
44519.4 50
0
9 Terminal~
194 741 598 0 1 3
0 31
0
0 0 49520 90
3 se1
-35 -6 -14 2
3 T44
-10 -32 11 -24
0
4 se1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3153 0 0
2
44519.4 51
0
9 Terminal~
194 741 589 0 1 3
0 29
0
0 0 49520 90
3 sn1
-35 -6 -14 2
3 T43
-10 -32 11 -24
0
4 sn1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
634 0 0
2
44519.4 52
0
9 Terminal~
194 741 580 0 1 3
0 31
0
0 0 49520 90
3 se2
-36 -5 -15 3
3 T42
-10 -32 11 -24
0
4 se2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8956 0 0
2
44519.4 53
0
9 Terminal~
194 741 571 0 1 3
0 27
0
0 0 49520 90
3 sn2
-35 -6 -14 2
3 T41
-10 -32 11 -24
0
4 sn2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3342 0 0
2
44519.4 54
0
9 Terminal~
194 741 562 0 1 3
0 31
0
0 0 49520 90
3 se3
-36 -6 -15 2
3 T40
-10 -32 11 -24
0
4 se3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3549 0 0
2
44519.4 55
0
9 Terminal~
194 741 553 0 1 3
0 26
0
0 0 49520 90
3 sn3
-35 -6 -14 2
3 T39
-10 -32 11 -24
0
4 sn3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9177 0 0
2
44519.4 56
0
7 Ground~
168 739 645 0 1 3
0 9
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3387 0 0
2
44519.4 57
0
7 74LS157
122 784 578 0 14 29
0 34 26 31 27 31 29 31 28 30
9 76 75 74 73
0
0 0 4848 0
7 74LS157
-24 -60 25 -52
2 U6
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
351 0 0
2
44519.4 58
0
7 Ground~
168 711 201 0 1 3
0 9
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3127 0 0
2
44519.4 59
0
9 Terminal~
194 600 196 0 1 3
0 30
0
0 0 49520 90
6 clock3
-50 -5 -8 3
3 T22
-10 -32 11 -24
0
7 clock3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
559 0 0
2
44519.4 60
0
9 Terminal~
194 600 205 0 1 3
0 25
0
0 0 49520 90
6 clock2
-49 -5 -7 3
3 T21
-10 -32 11 -24
0
7 clock2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8488 0 0
2
44519.4 61
0
9 Terminal~
194 600 169 0 1 3
0 35
0
0 0 49520 90
7 coluna3
-55 -7 -6 1
3 T20
-10 -32 11 -24
0
8 coluna3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3392 0 0
2
44519.4 62
0
9 Terminal~
194 600 178 0 1 3
0 36
0
0 0 49520 90
7 coluna2
-55 -7 -6 1
3 T19
-10 -32 11 -24
0
8 coluna2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3952 0 0
2
44519.4 63
0
9 Terminal~
194 600 187 0 1 3
0 37
0
0 0 49520 90
7 coluna1
-55 -7 -6 1
3 T18
-10 -32 11 -24
0
8 coluna1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8186 0 0
2
44519.4 64
0
9 Terminal~
194 514 366 0 1 3
0 35
0
0 0 49520 180
7 coluna3
4 -7 53 1
3 T17
-10 -32 11 -24
0
8 coluna3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6571 0 0
2
44519.4 65
0
9 Terminal~
194 433 368 0 1 3
0 36
0
0 0 49520 180
7 coluna2
4 -7 53 1
3 T16
-10 -32 11 -24
0
8 coluna2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6167 0 0
2
44519.4 66
0
9 Terminal~
194 343 367 0 1 3
0 37
0
0 0 49520 180
7 coluna1
4 -7 53 1
3 T15
-10 -32 11 -24
0
8 coluna1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3566 0 0
2
44519.4 67
0
7 74LS153
119 665 194 0 14 29
0 113 35 36 37 30 25 114 115 116
117 9 118 32 119
0
0 0 4848 0
7 74LS153
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 512 1 0 0 0
1 U
3371 0 0
2
44519.4 68
0
9 Terminal~
194 282 532 0 1 3
0 30
0
0 0 49520 270
6 clock3
2 -4 44 4
3 T14
-10 -32 11 -24
0
7 clock3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4395 0 0
2
44519.4 69
0
9 Terminal~
194 282 541 0 1 3
0 25
0
0 0 49520 270
6 clock2
2 -5 44 3
3 T13
-10 -32 11 -24
0
7 clock2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6822 0 0
2
44519.4 70
0
2 +V
167 343 55 0 1 3
0 77
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8953 0 0
2
44519.4 71
0
9 Terminal~
194 206 155 0 1 3
0 22
0
0 0 49520 90
6 linha1
-21 -15 21 -7
3 T12
-10 -32 11 -24
0
7 linha1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4635 0 0
2
44519.4 72
0
9 Terminal~
194 206 218 0 1 3
0 24
0
0 0 49520 90
6 linha2
-21 -15 21 -7
3 T11
-10 -32 11 -24
0
7 linha2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6596 0 0
2
44519.4 73
0
9 Terminal~
194 204 281 0 1 3
0 23
0
0 0 49520 90
6 linha3
-21 -15 21 -7
3 T10
-10 -32 11 -24
0
7 linha3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3813 0 0
2
44519.4 74
0
9 Terminal~
194 205 344 0 1 3
0 34
0
0 0 49520 90
6 linha4
-21 -15 21 -7
2 T9
-7 -32 7 -24
0
7 linha4;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5639 0 0
2
44519.4 75
0
9 Terminal~
194 233 646 0 1 3
0 24
0
0 0 49520 270
6 linha2
2 -5 44 3
2 T8
-7 -32 7 -24
0
7 linha2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
429 0 0
2
44519.4 76
0
9 Terminal~
194 233 655 0 1 3
0 22
0
0 0 49520 270
6 linha1
2 -4 44 4
2 T7
-7 -32 7 -24
0
7 linha1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5832 0 0
2
44519.4 77
0
9 Terminal~
194 233 637 0 1 3
0 23
0
0 0 49520 270
6 linha3
2 -4 44 4
2 T6
-7 -32 7 -24
0
7 linha3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8856 0 0
2
44519.4 78
0
9 Terminal~
194 233 628 0 1 3
0 34
0
0 0 49520 270
6 linha4
2 -4 44 4
2 T5
-7 -32 7 -24
0
7 linha4;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
469 0 0
2
44519.4 79
0
7 74LS139
118 181 654 0 14 29
0 39 38 9 120 121 122 34 23 24
22 123 124 125 126
0
0 0 4848 0
7 74LS139
-24 -51 25 -43
2 U3
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
113 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+[%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 13 14 15 7 6 5
4 9 10 11 12 3 2 1 13 14
15 7 6 5 4 9 10 11 12 0
65 0 0 512 1 0 0 0
1 U
4529 0 0
2
44519.4 80
0
9 Terminal~
194 98 647 0 1 3
0 38
0
0 0 49520 90
6 clock0
-48 -4 -6 4
2 T4
-7 -32 7 -24
0
7 clock0;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
88 0 0
2
44519.4 81
0
9 Terminal~
194 98 638 0 1 3
0 39
0
0 0 49520 90
6 clock1
-45 -6 -3 2
2 T3
-7 -32 7 -24
0
7 clock1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3894 0 0
2
44519.4 82
0
9 Terminal~
194 282 559 0 1 3
0 38
0
0 0 49520 270
6 clock0
2 -5 44 3
2 T2
-7 -32 7 -24
0
7 clock0;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6890 0 0
2
44519.4 83
0
9 Terminal~
194 282 550 0 1 3
0 39
0
0 0 49520 270
6 clock1
2 -4 44 4
2 T1
-7 -32 7 -24
0
7 clock1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3257 0 0
2
44519.4 84
0
7 Ground~
168 135 721 0 1 3
0 9
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6612 0 0
2
44519.4 85
0
7 74LS293
154 190 540 0 8 17
0 9 9 72 38 30 25 39 38
0
0 0 4848 0
7 74LS293
-24 -35 25 -27
2 U1
-7 -36 7 -28
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 0 1 0 0 0
1 U
3556 0 0
2
44519.4 86
0
7 Pulser~
4 74 474 0 10 12
0 127 128 5 40 0 0 10 10 3
7
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9143 0 0
2
44519.4 87
0
14 NO PushButton~
191 477 317 0 2 5
0 35 34
0
0 0 4208 0
0
3 S15
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
8186 0 0
2
44519.4 88
0
14 NO PushButton~
191 396 316 0 2 5
0 36 34
0
0 0 4208 0
0
3 S14
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3754 0 0
2
44519.4 89
0
14 NO PushButton~
191 314 316 0 2 5
0 37 34
0
0 0 4208 0
0
3 S13
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
8708 0 0
2
44519.4 90
0
14 NO PushButton~
191 478 254 0 2 5
0 35 23
0
0 0 4208 0
0
3 S11
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3338 0 0
2
44519.4 91
0
14 NO PushButton~
191 397 253 0 2 5
0 36 23
0
0 0 4208 0
0
3 S10
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
5546 0 0
2
44519.4 92
0
14 NO PushButton~
191 315 253 0 2 5
0 37 23
0
0 0 4208 0
0
2 S9
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3295 0 0
2
44519.4 93
0
14 NO PushButton~
191 478 191 0 2 5
0 35 24
0
0 0 4208 0
0
2 S7
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
4923 0 0
2
44519.4 94
0
14 NO PushButton~
191 397 190 0 2 5
0 36 24
0
0 0 4208 0
0
2 S5
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3248 0 0
2
44519.4 95
0
14 NO PushButton~
191 315 190 0 2 5
0 37 24
0
0 0 4208 0
0
2 S4
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3139 0 0
2
44519.4 96
0
14 NO PushButton~
191 477 128 0 2 5
0 35 22
0
0 0 4208 0
0
2 S3
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3285 0 0
2
44519.4 97
0
14 NO PushButton~
191 396 127 0 2 5
0 36 22
0
0 0 4208 0
0
2 S2
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
336 0 0
2
44519.4 98
0
14 NO PushButton~
191 314 127 0 2 5
0 37 22
0
0 0 4208 0
0
2 S1
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
6582 0 0
2
44519.4 99
0
9 Resistor~
219 433 90 0 4 5
0 36 77 0 1
0
0 0 880 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3546 0 0
2
44519.4 100
0
9 Resistor~
219 514 89 0 4 5
0 35 77 0 1
0
0 0 880 90
2 1k
8 0 22 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
893 0 0
2
44519.4 101
0
9 Resistor~
219 343 89 0 4 5
0 37 77 0 1
0
0 0 880 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8998 0 0
2
44519.4 102
0
205
4 1 40 0 0 4224 0 154 1 0 0 4
104 474
129 474
129 485
154 485
2 2 41 0 0 4224 0 9 13 0 0 2
1347 1504
1362 1504
3 1 2 0 0 4096 0 13 10 0 0 2
1407 1495
1438 1495
1 1 3 0 0 8192 0 11 9 0 0 3
1267 1502
1267 1504
1311 1504
1 1 4 0 0 4224 0 13 12 0 0 2
1362 1486
1304 1486
3 1 2 0 0 0 0 14 17 0 0 2
1103 1495
1134 1495
1 2 3 0 0 0 0 16 14 0 0 3
1035 1503
1035 1504
1058 1504
1 1 5 0 0 4224 0 14 15 0 0 2
1058 1486
1000 1486
1 1 9 0 0 12288 0 18 23 0 0 4
1710 1238
1710 1220
1681 1220
1681 1331
6 1 8 0 0 4224 0 18 22 0 0 3
1734 1259
1792 1259
1792 1258
1 4 7 0 0 4224 0 21 18 0 0 3
1642 1313
1710 1313
1710 1301
3 1 6 0 0 4224 0 18 20 0 0 3
1686 1277
1609 1277
1609 1275
1 2 42 0 0 8320 0 19 18 0 0 3
1649 1256
1649 1259
1686 1259
1 1 9 0 0 0 0 24 29 0 0 4
1400 1238
1400 1220
1371 1220
1371 1331
6 1 11 0 0 4224 0 24 28 0 0 3
1424 1259
1482 1259
1482 1258
1 4 10 0 0 4224 0 27 24 0 0 3
1332 1313
1400 1313
1400 1301
3 1 2 0 0 4224 0 24 26 0 0 3
1376 1277
1299 1277
1299 1275
1 2 43 0 0 8320 0 25 24 0 0 3
1339 1256
1339 1259
1376 1259
12 1 3 0 0 4224 0 41 30 0 0 2
1725 1042
1792 1042
1 1 9 0 0 0 0 36 31 0 0 4
1105 1239
1105 1221
1076 1221
1076 1332
6 1 12 0 0 4224 0 36 32 0 0 3
1129 1260
1187 1260
1187 1259
1 4 13 0 0 4224 0 33 36 0 0 3
1037 1314
1105 1314
1105 1302
3 1 14 0 0 4224 0 36 34 0 0 3
1081 1278
1004 1278
1004 1276
1 2 44 0 0 8320 0 35 36 0 0 3
1044 1257
1044 1260
1081 1260
3 1 45 0 0 8320 0 41 38 0 0 3
1655 1015
1620 1015
1620 951
8 0 9 0 0 0 0 41 0 0 29 2
1661 1060
1645 1060
7 0 9 0 0 0 0 41 0 0 29 2
1661 1051
1645 1051
6 0 9 0 0 0 0 41 0 0 29 2
1661 1042
1645 1042
5 1 9 0 0 0 0 41 37 0 0 3
1661 1033
1645 1033
1645 1111
0 4 9 0 0 0 0 0 41 29 0 3
1645 1033
1645 1024
1661 1024
1 2 15 0 0 8320 0 39 41 0 0 3
1600 1003
1600 1006
1661 1006
1 1 16 0 0 4224 0 41 40 0 0 2
1661 997
1639 997
1 1 17 0 0 4224 0 42 45 0 0 2
1342 998
1260 998
3 1 46 0 0 8320 0 42 44 0 0 3
1336 1016
1292 1016
1292 964
2 0 9 0 0 0 0 42 0 0 36 3
1342 1007
1326 1007
1326 1025
0 4 9 0 0 0 0 0 42 40 0 3
1326 1034
1326 1025
1342 1025
8 0 9 0 0 0 0 42 0 0 40 2
1342 1061
1325 1061
7 0 9 0 0 0 0 42 0 0 40 2
1342 1052
1325 1052
6 0 9 0 0 0 0 42 0 0 40 2
1342 1043
1325 1043
5 1 9 0 0 0 0 42 43 0 0 3
1342 1034
1325 1034
1325 1107
13 -207997 47 0 0 4224 0 63 0 0 45 2
1991 321
2062 321
14 -207998 48 0 0 4224 0 63 0 0 45 2
1991 330
2062 330
15 -207999 49 0 0 4224 0 63 0 0 45 2
1991 339
2062 339
16 -208000 50 0 0 4224 0 63 0 0 45 2
1991 348
2062 348
-13308169 0 1 0 0 4128 0 0 0 0 0 2
2062 138
2062 707
1 19 51 0 0 8320 0 2 65 0 0 4
1680 296
1724 296
1724 368
1710 368
18 0 52 0 0 12416 0 63 0 0 78 4
1991 276
2002 276
2002 217
1741 217
1 17 9 0 0 0 0 46 63 0 0 3
1904 296
1904 276
1921 276
5 -3261 53 0 0 4096 0 63 0 0 77 2
1927 321
1823 321
6 -3262 54 0 0 4096 0 63 0 0 77 2
1927 330
1823 330
7 -3263 55 0 0 4096 0 63 0 0 77 2
1927 339
1823 339
3 0 56 0 0 4096 0 47 0 0 55 2
2517 207
2435 207
3 0 56 0 0 0 0 54 0 0 55 2
2514 349
2435 349
3 0 56 0 0 0 0 58 0 0 55 2
2514 497
2435 497
1 3 56 0 0 8320 0 7 62 0 0 4
2422 149
2435 149
2435 637
2517 637
6 1 57 0 0 4224 0 62 59 0 0 2
2565 619
2611 619
4 1 9 0 0 0 0 62 60 0 0 2
2541 661
2541 673
1 1 9 0 0 0 0 62 61 0 0 4
2541 598
2541 559
2641 559
2641 572
1 2 58 0 0 4224 0 6 62 0 0 2
2487 619
2517 619
6 1 59 0 0 4224 0 58 55 0 0 2
2562 479
2608 479
4 1 9 0 0 0 0 58 56 0 0 2
2538 521
2538 533
1 1 9 0 0 0 0 58 57 0 0 4
2538 458
2538 419
2645 419
2645 428
1 2 60 0 0 4224 0 5 58 0 0 2
2484 479
2514 479
6 1 61 0 0 4224 0 54 51 0 0 2
2562 331
2610 331
4 1 9 0 0 0 0 54 52 0 0 2
2538 373
2538 387
1 1 9 0 0 0 0 54 53 0 0 4
2538 310
2538 273
2645 273
2645 284
1 2 62 0 0 4224 0 4 54 0 0 2
2482 331
2514 331
6 1 63 0 0 4224 0 47 50 0 0 2
2565 189
2611 189
4 1 9 0 0 0 0 47 49 0 0 2
2541 231
2541 243
1 1 9 0 0 0 0 47 48 0 0 4
2541 168
2541 129
2647 129
2647 143
1 2 64 0 0 4224 0 3 47 0 0 2
2487 189
2517 189
8 -3264 65 0 0 4096 0 63 0 0 77 2
1927 348
1823 348
15 -3261 53 0 0 4224 0 65 0 0 77 2
1704 422
1823 422
16 -3262 54 0 0 4224 0 65 0 0 77 2
1704 431
1823 431
17 -3263 55 0 0 4224 0 65 0 0 77 2
1704 440
1823 440
18 -3264 65 0 0 4224 0 65 0 0 77 2
1704 449
1823 449
-846037834 0 1 0 0 32 0 0 0 0 0 2
1823 140
1823 709
1 20 52 0 0 0 0 8 65 0 0 4
1608 154
1741 154
1741 377
1710 377
6 0 9 0 0 0 0 65 0 0 84 2
1640 413
1624 413
5 0 9 0 0 0 0 65 0 0 84 2
1640 404
1624 404
4 0 9 0 0 0 0 65 0 0 84 2
1640 395
1624 395
3 0 9 0 0 0 0 65 0 0 84 2
1640 386
1624 386
2 0 9 0 0 0 0 65 0 0 84 2
1640 377
1624 377
1 1 9 0 0 0 0 65 64 0 0 3
1640 368
1624 368
1624 473
7 -3453 66 0 0 4224 0 65 0 0 93 2
1640 422
1522 422
8 -3454 67 0 0 4224 0 65 0 0 93 2
1640 431
1522 431
9 -3455 68 0 0 4224 0 65 0 0 93 2
1640 440
1522 440
10 -3456 69 0 0 4224 0 65 0 0 93 2
1640 449
1522 449
4 -3453 66 0 0 0 0 66 0 0 93 3
1237 328
1237 436
1332 436
3 -3454 67 0 0 0 0 66 0 0 93 3
1243 328
1243 416
1332 416
2 -3455 68 0 0 0 0 66 0 0 93 3
1249 328
1249 401
1332 401
1 -3456 69 0 0 0 0 66 0 0 93 3
1255 328
1255 378
1332 378
-203315 0 1 0 0 12448 0 0 0 0 0 4
1332 728
1332 136
1522 136
1522 732
0 1 31 0 0 8192 0 0 92 117 0 3
555 721
555 730
572 730
2 1 70 0 0 4224 0 67 69 0 0 2
783 176
797 176
2 1 5 0 0 0 0 69 68 0 0 3
797 194
775 194
775 202
1 3 18 0 0 0 0 70 71 0 0 2
86 203
86 203
1 4 21 0 0 0 0 74 71 0 0 2
80 203
80 203
1 2 20 0 0 0 0 73 71 0 0 2
92 203
92 203
1 1 19 0 0 0 0 72 71 0 0 2
98 203
98 203
2 0 9 0 0 0 0 75 0 0 108 2
515 542
506 542
4 1 25 0 0 4096 0 75 81 0 0 2
515 560
494 560
1 3 30 0 0 4096 0 86 75 0 0 2
494 551
515 551
1 13 28 0 0 4224 0 84 75 0 0 2
604 587
579 587
1 12 29 0 0 4224 0 85 75 0 0 2
604 578
579 578
1 11 27 0 0 4224 0 83 75 0 0 2
604 569
579 569
1 10 26 0 0 4224 0 82 75 0 0 2
604 560
579 560
1 0 9 0 0 0 0 75 0 0 110 3
515 533
506 533
506 569
9 0 9 0 0 0 0 75 0 0 110 2
515 614
506 614
5 1 9 0 0 0 0 75 80 0 0 3
515 569
506 569
506 629
1 8 24 0 0 4096 0 79 75 0 0 2
500 596
515 596
2 7 71 0 0 4224 0 76 75 0 0 2
441 587
515 587
1 1 23 0 0 4096 0 78 76 0 0 2
404 587
405 587
1 6 22 0 0 4096 0 77 75 0 0 2
500 578
515 578
1 1 25 0 0 0 0 87 88 0 0 2
494 721
501 721
1 1 30 0 0 4096 0 91 93 0 0 2
572 739
546 739
1 2 31 0 0 4224 0 90 88 0 0 2
572 721
537 721
1 0 31 0 0 0 0 89 0 0 117 3
572 712
548 712
548 721
3 1 33 0 0 4096 0 69 111 0 0 2
842 185
860 185
0 1 5 0 0 0 0 0 94 122 0 2
117 465
154 465
3 3 72 0 0 4224 0 95 153 0 0 2
126 549
152 549
1 3 5 0 0 128 0 95 154 0 0 6
81 540
63 540
63 514
117 514
117 465
98 465
1 2 32 0 0 4096 0 96 95 0 0 2
69 558
81 558
0 1 32 0 0 8192 0 0 97 156 0 3
721 176
721 135
765 135
14 2 73 0 0 8320 0 125 98 0 0 4
816 614
873 614
873 711
950 711
13 2 74 0 0 4224 0 125 102 0 0 3
816 596
947 596
947 594
2 12 75 0 0 8320 0 106 125 0 0 4
944 483
873 483
873 578
816 578
11 2 76 0 0 8320 0 125 114 0 0 4
816 560
864 560
864 370
942 370
1 3 33 0 0 0 0 101 98 0 0 2
949 729
950 729
6 1 19 0 0 4224 0 98 100 0 0 2
998 711
1055 711
1 1 9 0 0 0 0 98 99 0 0 3
974 690
1026 690
1026 754
4 1 9 0 0 0 0 98 99 0 0 3
974 753
974 754
1026 754
1 3 33 0 0 0 0 105 102 0 0 2
932 612
947 612
6 1 20 0 0 4224 0 102 104 0 0 2
995 594
1052 594
1 1 9 0 0 0 0 102 103 0 0 3
971 573
1023 573
1023 637
4 1 9 0 0 0 0 102 103 0 0 3
971 636
971 637
1023 637
1 3 33 0 0 0 0 109 106 0 0 2
931 501
944 501
6 1 18 0 0 4224 0 106 108 0 0 2
992 483
1049 483
1 1 9 0 0 0 0 106 107 0 0 3
968 462
1020 462
1020 526
4 1 9 0 0 0 0 106 107 0 0 3
968 525
968 526
1020 526
1 3 33 0 0 4224 0 110 114 0 0 2
923 388
942 388
6 1 21 0 0 4224 0 114 112 0 0 2
990 370
1047 370
1 1 9 0 0 0 0 114 113 0 0 3
966 349
1018 349
1018 413
4 1 9 0 0 0 0 114 113 0 0 3
966 412
966 413
1018 413
1 1 34 0 0 0 0 115 125 0 0 2
752 542
752 542
1 8 28 0 0 0 0 117 125 0 0 2
752 605
752 605
1 9 30 0 0 0 0 116 125 0 0 2
752 614
752 614
1 6 29 0 0 0 0 119 125 0 0 4
752 587
753 587
753 587
752 587
1 7 31 0 0 0 0 118 125 0 0 2
752 596
752 596
1 4 27 0 0 0 0 121 125 0 0 2
752 569
752 569
1 5 31 0 0 0 0 120 125 0 0 2
752 578
752 578
1 2 26 0 0 0 0 123 125 0 0 2
752 551
752 551
1 3 31 0 0 0 0 122 125 0 0 2
752 560
752 560
1 10 9 0 0 0 0 124 125 0 0 3
739 639
739 623
746 623
1 11 9 0 0 0 0 126 135 0 0 3
711 195
711 158
703 158
13 1 32 0 0 4224 0 135 67 0 0 2
697 176
747 176
1 5 30 0 0 0 0 127 135 0 0 2
611 194
633 194
1 6 25 0 0 4096 0 128 135 0 0 2
611 203
633 203
1 2 35 0 0 4096 0 129 135 0 0 2
611 167
633 167
1 3 36 0 0 4096 0 130 135 0 0 2
611 176
633 176
1 4 37 0 0 4096 0 131 135 0 0 2
611 185
633 185
6 1 25 0 0 4224 0 153 137 0 0 2
222 540
270 540
5 1 30 0 0 4224 0 153 136 0 0 2
222 531
270 531
2 0 9 0 0 0 0 153 0 0 165 2
158 540
135 540
0 1 9 0 0 4224 0 0 153 200 0 3
135 654
135 531
158 531
2 0 22 0 0 4096 0 166 0 0 195 2
297 135
297 153
2 0 22 0 0 0 0 165 0 0 195 2
379 135
379 153
2 0 24 0 0 4096 0 163 0 0 194 2
298 198
298 216
2 0 24 0 0 0 0 162 0 0 194 2
380 198
380 216
2 0 23 0 0 4096 0 160 0 0 193 2
298 261
298 279
2 0 23 0 0 0 0 159 0 0 193 2
380 261
380 279
2 0 34 0 0 4096 0 157 0 0 192 2
297 324
297 342
2 0 34 0 0 0 0 156 0 0 192 2
379 324
379 342
1 0 35 0 0 0 0 155 0 0 188 2
494 325
514 325
1 0 35 0 0 0 0 158 0 0 188 2
495 262
514 262
1 0 35 0 0 0 0 161 0 0 188 2
495 199
514 199
1 0 36 0 0 0 0 156 0 0 189 2
413 324
433 324
1 0 36 0 0 0 0 159 0 0 189 2
414 261
433 261
1 0 36 0 0 0 0 162 0 0 189 2
414 198
433 198
1 0 37 0 0 0 0 157 0 0 190 2
331 324
343 324
1 0 37 0 0 0 0 160 0 0 190 2
332 261
343 261
1 0 37 0 0 0 0 163 0 0 190 2
332 198
343 198
1 0 35 0 0 0 0 164 0 0 188 2
494 136
514 136
1 0 36 0 0 0 0 165 0 0 189 2
413 135
433 135
1 0 37 0 0 0 0 166 0 0 190 2
331 135
343 135
2 2 77 0 0 8192 0 167 168 0 0 3
433 72
433 71
514 71
2 2 77 0 0 4224 0 169 167 0 0 3
343 71
433 71
433 72
1 1 35 0 0 4224 0 168 132 0 0 2
514 107
514 351
1 1 36 0 0 4224 0 167 133 0 0 2
433 108
433 353
1 1 37 0 0 4224 0 169 134 0 0 2
343 107
343 352
2 1 77 0 0 0 0 169 138 0 0 2
343 71
343 64
1 2 34 0 0 4224 0 142 155 0 0 3
216 342
460 342
460 325
1 2 23 0 0 4224 0 141 158 0 0 3
215 279
461 279
461 262
1 2 24 0 0 4224 0 140 161 0 0 3
217 216
461 216
461 199
1 2 22 0 0 4224 0 139 164 0 0 3
217 153
460 153
460 136
1 10 22 0 0 0 0 144 147 0 0 2
221 654
219 654
1 9 24 0 0 0 0 143 147 0 0 2
221 645
219 645
1 8 23 0 0 0 0 145 147 0 0 2
221 636
219 636
1 7 34 0 0 0 0 146 147 0 0 2
221 627
219 627
3 1 9 0 0 0 0 147 152 0 0 3
143 654
135 654
135 715
1 2 38 0 0 4096 0 148 147 0 0 2
109 645
149 645
1 1 39 0 0 4096 0 149 147 0 0 2
109 636
149 636
0 1 38 0 0 0 0 0 150 205 0 2
234 558
270 558
7 1 39 0 0 4224 0 153 151 0 0 2
222 549
270 549
8 4 38 0 0 12416 0 153 153 0 0 6
222 558
234 558
234 575
144 575
144 558
152 558
29
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 27
1318 1522 1453 1566
1325 1527 1445 1559
27 clock AND q!=4:
   or_down
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 24
1016 1521 1143 1565
1023 1526 1135 1558
24 clock AND q=4:
   or_up
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
1720 1325 1823 1349
1727 1330 1815 1346
11 ddisponivel
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1401 1323 1472 1347
1408 1329 1464 1345
7 overrun
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1101 1319 1156 1343
1108 1324 1148 1340
5 write
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
1646 1082 1741 1106
1653 1087 1733 1103
10 quantidade
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1342 1080 1405 1104
1349 1086 1397 1102
6 inicio
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 41
917 162 1096 206
922 166 1090 198
41 set ao clicar o botao
e ao subir o clock
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
64 73 119 97
71 78 111 94
5 saida
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
1143 507 1226 551
1148 511 1220 543
20 "memoria"
de 4 bits
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 51
675 450 838 514
680 454 832 502
51 multiplex para
escolher entre
as duas aritmeticas
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 24
437 672 640 696
442 676 634 692
24 aritmetica para *, 0 e #
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
454 479 617 503
459 483 611 499
19 aritmetica para 1-9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
147 428 282 452
150 430 278 446
16 divisao do clock
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
299 288 330 312
302 290 326 306
3 (*)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
462 289 493 313
465 291 489 307
3 (#)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
381 288 412 312
384 290 408 306
3 (0)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
463 226 494 250
466 228 490 244
3 (9)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
382 225 413 249
385 227 409 243
3 (8)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
300 225 331 249
303 227 327 243
3 (7)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
463 163 494 187
466 165 490 181
3 (6)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
382 162 413 186
385 164 409 180
3 (5)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
300 162 331 186
303 164 327 180
3 (4)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
462 99 493 123
465 101 489 117
3 (3)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
381 98 412 122
384 100 408 116
3 (2)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
295 93 334 117
302 99 326 115
3 (1)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
397 37 540 61
404 42 532 58
16 matriz de botoes
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
55 93 120 132
63 100 111 130
14 * -> E
# -> F
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 82
2353 60 2736 102
2365 70 2723 100
82 REGISTRADOR (Entradas tempor�rias com chaves s� pra 
mostrar que t� funcionando)
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
