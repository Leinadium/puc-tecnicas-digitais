CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
1140 910 2 120 10
176 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.331203 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
234
13 Logic Switch~
5 1936 1350 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9154 0 0
2
44519.9 0
0
13 Logic Switch~
5 1560 965 0 10 11
0 51 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V13
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8600 0 0
2
44519.9 0
0
13 Logic Switch~
5 2475 189 0 1 11
0 86
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6288 0 0
2
44519.9 1
0
13 Logic Switch~
5 2470 331 0 1 11
0 84
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5914 0 0
2
44519.9 2
0
13 Logic Switch~
5 2472 479 0 1 11
0 82
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9916 0 0
2
44519.9 3
0
13 Logic Switch~
5 2475 619 0 1 11
0 80
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
946 0 0
2
44519.9 4
0
13 Logic Switch~
5 2410 149 0 1 11
0 78
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7876 0 0
2
44519.9 5
0
13 Logic Switch~
5 1596 154 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4411 0 0
2
44519.9 6
0
7 Ground~
168 1679 1321 0 1 3
0 2
0
0 0 53360 0
0
5 GND20
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
836 0 0
2
44519.9 0
0
2 +V
167 1663 1235 0 1 3
0 49
0
0 0 54256 0
2 5V
-7 -22 7 -14
3 V11
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3878 0 0
2
44519.9 0
0
9 Terminal~
194 1710 1328 0 1 3
0 3
0
0 0 49520 180
6 dddown
7 -7 49 1
3 T65
-11 -32 10 -24
0
7 dddown;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4956 0 0
2
44519.9 0
0
14 Logic Display~
6 1843 1244 0 1 2
10 28
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3765 0 0
2
44519.9 0
0
9 Terminal~
194 1973 1343 0 1 3
0 4
0
0 0 49520 0
4 wrup
-14 -22 14 -14
3 T89
-11 -32 10 -24
0
5 wrup;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7205 0 0
2
44519.9 1
0
2 +V
167 1293 946 0 1 3
0 50
0
0 0 54256 0
2 5V
-7 -22 7 -14
3 V10
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4258 0 0
2
44519.9 0
0
9 Terminal~
194 1177 1616 0 1 3
0 5
0
0 0 49520 0
2 pq
-7 -22 7 -14
4 T115
-14 -32 14 -24
0
3 pq;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5549 0 0
2
44519.9 0
0
7 74LS191
135 1641 1024 0 14 29
0 2 5 51 10 2 2 2 2 95
96 9 6 7 8
0
0 0 4848 0
7 74LS191
-24 -51 25 -43
3 U25
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 0 0 0 0
1 U
6519 0 0
2
44519.9 8
0
9 Terminal~
194 1699 1043 0 1 3
0 6
0
0 0 49520 270
4 qua3
6 -7 34 1
4 T130
-13 -32 15 -24
0
5 qua3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6340 0 0
2
44519.9 7
0
9 Terminal~
194 1699 1052 0 1 3
0 7
0
0 0 49520 270
4 qua2
6 -7 34 1
4 T131
-13 -32 15 -24
0
5 qua2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3158 0 0
2
44519.9 6
0
9 Terminal~
194 1699 1061 0 1 3
0 8
0
0 0 49520 270
4 qua1
5 -6 33 2
4 T132
-13 -32 15 -24
0
5 qua1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9342 0 0
2
44519.9 5
0
9 Terminal~
194 1739 1024 0 1 3
0 9
0
0 0 49520 0
5 qoito
-17 -22 18 -14
4 T133
-14 -32 14 -24
0
6 qoito;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8937 0 0
2
44519.9 4
0
7 Ground~
168 1592 1117 0 1 3
0 2
0
0 0 53360 0
0
5 GND24
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4688 0 0
2
44519.9 3
0
9 Terminal~
194 1567 1026 0 1 3
0 10
0
0 0 49520 90
4 modo
-35 -6 -7 2
4 T134
-14 -32 14 -24
0
5 modo;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3401 0 0
2
44519.9 2
0
9 Terminal~
194 1567 1008 0 1 3
0 5
0
0 0 49520 90
2 pq
-28 -5 -14 3
4 T135
-14 -32 14 -24
0
3 pq;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4445 0 0
2
44519.9 1
0
9 Inverter~
13 1669 297 0 2 22
0 4 52
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 11 0
1 U
5487 0 0
2
44519.9 0
0
9 Terminal~
194 1619 288 0 1 3
0 4
0
0 0 49520 0
4 wrup
-14 -22 14 -14
4 T129
-14 -32 14 -24
0
5 wrup;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9241 0 0
2
44519.9 0
0
12 Hex Display~
7 1687 697 0 16 19
10 8 7 6 97 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 0 0 0 0
4 DISP
7598 0 0
2
44519.9 3
0
9 Terminal~
194 1684 761 0 1 3
0 6
0
0 0 49520 180
4 qua3
7 -7 35 1
4 T128
-13 -32 15 -24
0
5 qua3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7456 0 0
2
44519.9 2
0
9 Terminal~
194 1690 748 0 1 3
0 7
0
0 0 49520 180
4 qua2
7 -7 35 1
4 T127
-13 -32 15 -24
0
5 qua2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4625 0 0
2
44519.9 1
0
9 Terminal~
194 1696 736 0 1 3
0 8
0
0 0 49520 180
4 qua1
7 -7 35 1
4 T126
-13 -32 15 -24
0
5 qua1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9637 0 0
2
44519.9 0
0
9 Terminal~
194 1612 738 0 1 3
0 11
0
0 0 49520 180
4 ini1
7 -7 35 1
4 T124
-13 -32 15 -24
0
5 ini1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3175 0 0
2
44519.9 2
0
9 Terminal~
194 1606 750 0 1 3
0 12
0
0 0 49520 180
4 ini2
7 -7 35 1
3 T88
-10 -32 11 -24
0
5 ini2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4411 0 0
2
44519.9 1
0
9 Terminal~
194 1600 763 0 1 3
0 13
0
0 0 49520 180
4 ini3
7 -7 35 1
3 T87
-10 -32 11 -24
0
5 ini3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8285 0 0
2
44519.9 0
0
12 Hex Display~
7 1603 699 0 18 19
10 11 12 13 98 0 0 0 0 0
0 0 1 1 0 0 1 1 4
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 0 0 0 0
4 DISP
6178 0 0
2
44519.9 0
0
9 Terminal~
194 1774 155 0 1 3
0 10
0
0 0 49520 270
4 modo
6 -5 34 3
4 T104
-13 -32 15 -24
0
5 modo;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9911 0 0
2
44519.9 0
0
8 Hex Key~
166 2145 344 0 11 12
0 53 54 55 56 0 0 0 0 0
3 51
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
7251 0 0
2
44519.9 0
0
9 Terminal~
194 1623 1547 0 1 3
0 6
0
0 0 49520 90
4 qua3
-37 -6 -9 2
4 T118
-14 -32 14 -24
0
5 qua3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9851 0 0
2
44519.9 3
0
9 Terminal~
194 1623 1556 0 1 3
0 7
0
0 0 49520 90
4 qua2
-37 -6 -9 2
4 T119
-14 -32 14 -24
0
5 qua2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9133 0 0
2
44519.9 2
0
9 Terminal~
194 1623 1565 0 1 3
0 8
0
0 0 49520 90
4 qua1
-37 -6 -9 2
4 T120
-14 -32 14 -24
0
5 qua1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7576 0 0
2
44519.9 1
0
8 3-In OR~
219 1664 1554 0 4 22
0 6 7 8 57
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U24A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 14 0
1 U
9978 0 0
2
44519.9 0
0
9 Terminal~
194 1678 1460 0 1 3
0 10
0
0 0 49520 90
4 modo
-38 -6 -10 2
3 T84
-11 -32 10 -24
0
5 modo;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
758 0 0
2
44519.9 6
0
9 2-In AND~
219 1736 1467 0 3 22
0 10 14 3
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U23A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
5351 0 0
2
44519.9 5
0
9 Terminal~
194 1679 1478 0 1 3
0 14
0
0 0 49520 90
5 wrout
-41 -6 -6 2
4 T122
-14 -32 14 -24
0
6 wrout;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7860 0 0
2
44519.9 4
0
9 Terminal~
194 1807 1468 0 1 3
0 3
0
0 0 49520 270
6 dddown
-21 -15 21 -7
4 T123
-14 -32 14 -24
0
7 dddown;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8118 0 0
2
44519.9 3
0
9 Terminal~
194 1808 1524 0 1 3
0 15
0
0 0 49520 270
4 ddup
-15 -15 13 -7
4 T121
-14 -32 14 -24
0
5 ddup;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7363 0 0
2
44519.9 2
0
9 2-In AND~
219 1737 1523 0 3 22
0 16 57 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U23B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 13 0
1 U
9572 0 0
2
44519.9 1
0
9 Terminal~
194 1679 1516 0 1 3
0 16
0
0 0 49520 90
5 clock
-42 -6 -7 2
4 T125
-14 -32 14 -24
0
6 clock;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3608 0 0
2
44519.9 0
0
9 Terminal~
194 1294 746 0 1 3
0 9
0
0 0 49520 180
5 qoito
-13 11 22 19
3 T90
-10 -32 11 -24
0
6 qoito;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8671 0 0
2
44519.9 3
0
9 Terminal~
194 1276 745 0 1 3
0 6
0
0 0 49520 180
4 qua3
-20 1 8 9
3 T86
-10 -32 11 -24
0
5 qua3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9832 0 0
2
44519.9 2
0
8 2-In OR~
219 1282 695 0 3 22
0 6 9 60
0
0 0 624 90
6 74LS32
-21 -24 21 -16
4 U19C
29 -3 57 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
3630 0 0
2
44519.9 1
0
9 2-In AND~
219 1277 628 0 3 22
0 59 60 58
0
0 0 624 90
6 74LS08
-21 -24 21 -16
4 U20D
17 -5 45 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 10 0
1 U
3159 0 0
2
44519.9 0
0
9 Inverter~
13 1411 962 0 2 22
0 62 61
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U3B
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 11 0
1 U
7384 0 0
2
44519.9 0
0
9 Terminal~
194 1232 1674 0 1 3
0 17
0
0 0 49520 270
7 pinicio
-25 -15 24 -7
3 T85
-11 -32 10 -24
0
8 pinicio;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3933 0 0
2
44519.9 0
0
9 Terminal~
194 1036 1684 0 1 3
0 10
0
0 0 49520 90
4 modo
-36 -6 -8 2
4 T105
-14 -32 14 -24
0
5 modo;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8168 0 0
2
44519.9 0
0
5 4081~
219 1147 1673 0 3 22
0 5 10 17
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U22B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 12 0
1 U
5374 0 0
2
44519.9 0
0
9 Terminal~
194 1034 1618 0 1 3
0 14
0
0 0 49520 90
5 wrout
-39 -6 -4 2
4 T112
-14 -32 14 -24
0
6 wrout;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7500 0 0
2
44519.9 0
0
5 4081~
219 1085 1625 0 3 22
0 14 18 5
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U22A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 12 0
1 U
4207 0 0
2
44519.9 0
0
9 Terminal~
194 1130 1616 0 1 3
0 5
0
0 0 49520 0
6 wrdown
-21 -22 21 -14
4 T114
-14 -32 14 -24
0
7 wrdown;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3844 0 0
2
44519.9 0
0
9 Terminal~
194 1034 1636 0 1 3
0 18
0
0 0 49520 90
6 nclock
-43 -5 -1 3
4 T113
-14 -32 14 -24
0
7 nclock;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5174 0 0
2
44519.9 0
0
9 Terminal~
194 233 664 0 1 3
0 19
0
0 0 49520 270
7 clinha4
3 -4 52 4
4 T111
-14 -32 14 -24
0
8 clinha4;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5620 0 0
2
44519.9 7
0
9 Terminal~
194 233 673 0 1 3
0 20
0
0 0 49520 270
7 clinha3
1 -4 50 4
4 T110
-14 -32 14 -24
0
8 clinha3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5464 0 0
2
44519.9 8
0
9 Terminal~
194 233 691 0 1 3
0 21
0
0 0 49520 270
7 clinha1
2 -4 51 4
4 T109
-14 -32 14 -24
0
8 clinha1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5444 0 0
2
44519.9 9
0
9 Terminal~
194 233 682 0 1 3
0 22
0
0 0 49520 270
7 clinha2
2 -4 51 4
4 T108
-14 -32 14 -24
0
8 clinha2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3975 0 0
2
44519.9 10
0
9 Terminal~
194 96 674 0 1 3
0 23
0
0 0 49520 90
6 clock1
-45 -6 -3 2
4 T107
-14 -32 14 -24
0
7 clock1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5865 0 0
2
44519.9 11
0
9 Terminal~
194 96 683 0 1 3
0 24
0
0 0 49520 90
6 clock0
-48 -4 -6 4
4 T106
-14 -32 14 -24
0
7 clock0;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
859 0 0
2
44519.9 12
0
9 Terminal~
194 773 195 0 1 3
0 16
0
0 0 49520 90
5 clock
-45 -6 -10 2
3 T64
-10 -32 11 -24
0
6 clock;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4289 0 0
2
44519.9 17
0
9 2-In AND~
219 833 184 0 3 22
0 63 16 25
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U20C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 10 0
1 U
4623 0 0
2
44519.9 18
0
2 +V
167 617 127 0 1 3
0 64
0
0 0 54256 0
2 5V
-7 -22 7 -14
3 V12
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9733 0 0
2
44519.9 23
0
7 74LS139
118 181 654 0 14 29
0 23 24 2 23 24 2 42 48 47
46 19 20 22 21
0
0 0 13040 0
7 74LS139
-24 -51 25 -43
3 U21
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
113 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+[%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
13 type: digital
5 DIP16
29

0 3 2 1 13 14 15 7 6 5
4 9 10 11 12 3 2 1 13 14
15 7 6 5 4 9 10 11 12 70
65 0 0 0 1 1 0 0
1 U
4682 0 0
2
44519.9 24
0
7 74LS293
154 191 540 0 8 17
0 2 2 89 24 39 34 23 24
0
0 0 4848 0
7 74LS293
-24 -35 25 -27
2 U1
-7 -36 7 -28
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 0 1 0 0 0
1 U
8941 0 0
2
44519.9 25
0
9 Terminal~
194 918 185 0 1 3
0 25
0
0 0 49520 270
3 set
-17 6 4 14
3 T50
-10 -32 11 -24
0
4 set;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3820 0 0
2
5.90009e-315 0
0
9 Terminal~
194 1164 658 0 1 3
0 10
0
0 0 49520 90
4 modo
-32 -6 -4 2
3 T92
-10 -32 11 -24
0
5 modo;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8459 0 0
2
5.90009e-315 5.26354e-315
0
8 2-In OR~
219 1346 694 0 3 22
0 7 9 69
0
0 0 624 90
6 74LS32
-21 -24 21 -16
4 U19A
29 -3 57 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
3440 0 0
2
5.90009e-315 5.30499e-315
0
9 2-In AND~
219 1341 628 0 3 22
0 59 69 70
0
0 0 624 90
6 74LS08
-21 -24 21 -16
4 U20A
17 -5 45 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
5821 0 0
2
5.90009e-315 5.32571e-315
0
9 Inverter~
13 1221 656 0 2 22
0 10 59
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
775 0 0
2
5.90009e-315 5.34643e-315
0
9 Terminal~
194 1340 741 0 1 3
0 7
0
0 0 49520 180
4 qua2
-20 1 8 9
3 T91
-10 -32 11 -24
0
5 qua2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8472 0 0
2
5.90009e-315 5.3568e-315
0
9 Terminal~
194 1358 741 0 1 3
0 9
0
0 0 49520 180
5 qoito
-12 11 23 19
3 T93
-10 -32 11 -24
0
6 qoito;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5642 0 0
2
5.90009e-315 5.36716e-315
0
9 2-In AND~
219 1413 630 0 3 22
0 59 68 71
0
0 0 624 90
6 74LS08
-21 -24 21 -16
4 U20B
17 -5 45 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
5711 0 0
2
5.90009e-315 5.37752e-315
0
8 2-In OR~
219 1418 696 0 3 22
0 8 9 68
0
0 0 624 90
6 74LS32
-21 -24 21 -16
4 U19B
29 -3 57 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
8118 0 0
2
5.90009e-315 5.38788e-315
0
9 Terminal~
194 1412 743 0 1 3
0 8
0
0 0 49520 180
4 qua1
-20 1 8 9
3 T95
-10 -32 11 -24
0
5 qua1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3757 0 0
2
5.90009e-315 5.39306e-315
0
9 Terminal~
194 1430 743 0 1 3
0 9
0
0 0 49520 180
5 qoito
-13 11 22 19
4 T103
-13 -32 15 -24
0
6 qoito;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3882 0 0
2
5.90009e-315 5.39824e-315
0
9 Terminal~
194 1431 1044 0 1 3
0 13
0
0 0 49520 270
4 ini3
6 -6 34 2
3 T98
-10 -32 11 -24
0
5 ini3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9366 0 0
2
5.90009e-315 5.41378e-315
0
9 Terminal~
194 1431 1053 0 1 3
0 12
0
0 0 49520 270
4 ini2
6 -7 34 1
3 T99
-10 -32 11 -24
0
5 ini2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5650 0 0
2
5.90009e-315 5.41896e-315
0
9 Terminal~
194 1431 1062 0 1 3
0 11
0
0 0 49520 270
4 ini1
5 -6 33 2
4 T100
-13 -32 15 -24
0
5 ini1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7718 0 0
2
5.90009e-315 5.42414e-315
0
9 Terminal~
194 1447 523 0 1 3
0 13
0
0 0 49520 90
4 ini3
-32 -6 -4 2
3 T97
-10 -32 11 -24
0
5 ini3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6825 0 0
2
5.90009e-315 5.42933e-315
0
9 Terminal~
194 1447 532 0 1 3
0 12
0
0 0 49520 90
4 ini2
-32 -6 -4 2
3 T96
-10 -32 11 -24
0
5 ini2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8223 0 0
2
5.90009e-315 5.43192e-315
0
9 Terminal~
194 1447 541 0 1 3
0 11
0
0 0 49520 90
4 ini1
-32 -6 -4 2
3 T94
-10 -32 11 -24
0
5 ini1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4773 0 0
2
5.90009e-315 5.43451e-315
0
6 74LS83
105 1523 548 0 14 29
0 2 13 12 11 2 58 70 71 2
99 67 66 65 2
0
0 0 4848 0
6 74LS83
-21 -60 21 -52
3 U16
-10 -61 11 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
7329 0 0
2
5.90009e-315 5.4371e-315
0
7 Ground~
168 1475 664 0 1 3
0 2
0
0 0 53360 0
0
5 GND25
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5290 0 0
2
5.90009e-315 5.43969e-315
0
9 2-In AND~
219 1082 1495 0 3 22
0 16 9 27
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
6210 0 0
2
5.90009e-315 5.44228e-315
0
9 2-In AND~
219 1387 1495 0 3 22
0 18 72 26
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
4522 0 0
2
5.90009e-315 5.44487e-315
0
9 Terminal~
194 166 486 0 1 3
0 18
0
0 0 49520 270
6 nclock
2 -4 44 4
3 T83
-10 -32 11 -24
0
7 nclock;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4399 0 0
2
5.90009e-315 5.46818e-315
0
9 Inverter~
13 1326 1504 0 2 22
0 9 72
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
6836 0 0
2
5.90009e-315 5.47077e-315
0
9 Terminal~
194 1452 1486 0 1 3
0 26
0
0 0 49520 0
6 ordown
-21 -22 21 -14
3 T82
-11 -32 10 -24
0
7 ordown;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5657 0 0
2
5.90009e-315 5.47207e-315
0
9 Terminal~
194 1267 1493 0 1 3
0 9
0
0 0 49520 0
5 qoito
-17 -22 18 -14
3 T81
-11 -32 10 -24
0
6 qoito;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3900 0 0
2
5.90009e-315 5.47336e-315
0
9 Terminal~
194 1304 1477 0 1 3
0 18
0
0 0 49520 0
6 nclock
-20 -22 22 -14
3 T80
-11 -32 10 -24
0
7 nclock;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9532 0 0
2
5.90009e-315 5.47466e-315
0
9 Terminal~
194 1000 1477 0 1 3
0 16
0
0 0 49520 0
5 clock
-17 -22 18 -14
3 T77
-11 -32 10 -24
0
6 clock;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
347 0 0
2
5.90009e-315 5.47595e-315
0
9 Terminal~
194 1035 1494 0 1 3
0 9
0
0 0 49520 0
5 qoito
-17 -22 18 -14
3 T78
-11 -32 10 -24
0
6 qoito;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8304 0 0
2
5.90009e-315 5.47725e-315
0
9 Terminal~
194 1134 1486 0 1 3
0 27
0
0 0 49520 0
4 orup
-14 -22 14 -14
3 T79
-11 -32 10 -24
0
5 orup;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3414 0 0
2
5.90009e-315 5.47854e-315
0
5 4013~
219 1710 1295 0 6 22
0 2 49 15 3 100 28
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U18B
21 -54 49 -46
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 9 0
1 U
4979 0 0
2
5.90009e-315 5.47984e-315
0
9 Terminal~
194 1644 1267 0 1 3
0 15
0
0 0 49520 0
4 ddup
-14 -21 14 -13
3 T71
-11 -32 10 -24
0
5 ddup;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4312 0 0
2
5.90009e-315 5.48372e-315
0
9 Terminal~
194 1792 1249 0 1 3
0 28
0
0 0 49520 0
5 ddout
-17 -22 18 -14
3 T70
-11 -32 10 -24
0
6 ddout;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8210 0 0
2
5.90009e-315 5.48502e-315
0
5 4013~
219 1400 1295 0 6 22
0 2 73 27 26 101 29
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U18A
21 -54 49 -46
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 9 0
1 U
8709 0 0
2
5.90009e-315 5.48761e-315
0
2 +V
167 1339 1247 0 1 3
0 73
0
0 0 54256 0
3 10V
-11 -22 10 -14
3 V17
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8410 0 0
2
5.90009e-315 5.4889e-315
0
9 Terminal~
194 1299 1266 0 1 3
0 27
0
0 0 49520 0
4 orup
-14 -22 14 -14
3 T69
-11 -32 10 -24
0
5 orup;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6112 0 0
2
5.90009e-315 5.4902e-315
0
9 Terminal~
194 1332 1304 0 1 3
0 26
0
0 0 49520 0
6 ordown
-21 -22 21 -14
3 T68
-11 -32 10 -24
0
7 ordown;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4562 0 0
2
5.90009e-315 5.49149e-315
0
9 Terminal~
194 1482 1249 0 1 3
0 29
0
0 0 49520 0
5 orout
-17 -22 18 -14
3 T67
-11 -32 10 -24
0
6 orout;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3901 0 0
2
5.90009e-315 5.49279e-315
0
7 Ground~
168 1371 1337 0 1 3
0 2
0
0 0 53360 0
0
5 GND21
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5761 0 0
2
5.90009e-315 5.49408e-315
0
7 Ground~
168 1076 1338 0 1 3
0 2
0
0 0 53360 0
0
5 GND23
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
510 0 0
2
5.90009e-315 5.49667e-315
0
9 Terminal~
194 1187 1250 0 1 3
0 14
0
0 0 49520 0
5 wrout
-17 -22 18 -14
3 T75
-11 -32 10 -24
0
6 wrout;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3190 0 0
2
5.90009e-315 5.49797e-315
0
9 Terminal~
194 1037 1305 0 1 3
0 5
0
0 0 49520 0
6 wrdown
-21 -22 21 -14
3 T74
-11 -32 10 -24
0
7 wrdown;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
514 0 0
2
5.90009e-315 5.49926e-315
0
9 Terminal~
194 1004 1267 0 1 3
0 4
0
0 0 49520 0
4 wrup
-14 -22 14 -14
3 T73
-11 -32 10 -24
0
5 wrup;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7400 0 0
2
5.90009e-315 5.50056e-315
0
2 +V
167 1044 1248 0 1 3
0 74
0
0 0 54256 0
3 10V
-11 -22 10 -14
3 V16
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8722 0 0
2
5.90009e-315 5.50185e-315
0
5 4013~
219 1105 1296 0 6 22
0 2 74 4 5 102 14
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U17B
21 -54 49 -46
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 8 0
1 U
5565 0 0
2
5.90009e-315 5.50315e-315
0
7 74LS193
137 1374 1025 0 14 29
0 17 50 61 2 2 2 2 2 103
104 62 13 12 11
0
0 0 4848 0
7 74LS193
-24 -51 25 -43
3 U14
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
4511 0 0
2
5.90009e-315 5.51092e-315
0
7 Ground~
168 1325 1113 0 1 3
0 2
0
0 0 53360 0
0
5 GND19
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6586 0 0
2
5.90009e-315 5.51222e-315
0
9 Terminal~
194 1260 989 0 1 3
0 17
0
0 0 49520 0
7 pinicio
-25 -22 24 -14
3 T63
-11 -32 10 -24
0
8 pinicio;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8917 0 0
2
5.90009e-315 5.51351e-315
0
7 Ground~
168 1904 302 0 1 3
0 2
0
0 0 53360 0
0
5 GND18
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7921 0 0
2
44519.9 26
0
5 4013~
219 2541 225 0 6 22
0 2 86 78 2 105 85
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U10A
23 -61 51 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 5 0
1 U
6731 0 0
2
44519.9 27
0
7 Ground~
168 2647 149 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9825 0 0
2
44519.9 28
0
7 Ground~
168 2541 249 0 1 3
0 2
0
0 0 53360 0
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8689 0 0
2
44519.9 29
0
14 Logic Display~
6 2611 171 0 1 2
10 85
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
356 0 0
2
44519.9 30
0
14 Logic Display~
6 2610 313 0 1 2
10 83
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9622 0 0
2
44519.9 31
0
7 Ground~
168 2538 393 0 1 3
0 2
0
0 0 53360 0
0
5 GND11
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9335 0 0
2
44519.9 32
0
7 Ground~
168 2645 290 0 1 3
0 2
0
0 0 53360 0
0
5 GND12
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3748 0 0
2
44519.9 33
0
5 4013~
219 2538 367 0 6 22
0 2 84 78 2 106 83
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U10B
23 -61 51 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 5 0
1 U
8642 0 0
2
44519.9 34
0
14 Logic Display~
6 2608 461 0 1 2
10 81
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3377 0 0
2
44519.9 35
0
7 Ground~
168 2538 539 0 1 3
0 2
0
0 0 53360 0
0
5 GND13
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9599 0 0
2
44519.9 36
0
7 Ground~
168 2645 434 0 1 3
0 2
0
0 0 53360 0
0
5 GND14
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3104 0 0
2
44519.9 37
0
5 4013~
219 2538 515 0 6 22
0 2 82 78 2 107 81
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U11A
23 -61 51 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 6 0
1 U
3441 0 0
2
44519.9 38
0
14 Logic Display~
6 2611 601 0 1 2
10 79
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9765 0 0
2
44519.9 39
0
7 Ground~
168 2541 679 0 1 3
0 2
0
0 0 53360 0
0
5 GND15
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3229 0 0
2
44519.9 40
0
7 Ground~
168 2641 578 0 1 3
0 2
0
0 0 53360 0
0
5 GND16
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4643 0 0
2
44519.9 41
0
5 4013~
219 2541 655 0 6 22
0 2 80 78 2 108 79
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U11B
23 -61 51 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 6 0
1 U
4404 0 0
2
44519.9 42
0
7 74LS245
64 1959 312 0 18 37
0 109 110 111 112 75 76 77 87 113
114 115 116 56 55 54 53 2 10
0
0 0 4848 0
7 74LS245
-24 -60 25 -52
3 U13
-11 -61 10 -53
0
16 DVCC=20;DGND=10;
192 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i]
+ [%20bi %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP14
37

0 9 8 7 6 5 4 3 2 11
12 13 14 15 16 17 18 19 1 9
8 7 6 5 4 3 2 11 12 13
14 15 16 17 18 19 1 0
65 0 0 512 1 0 0 0
1 U
5170 0 0
2
44519.9 43
0
7 Ground~
168 1624 479 0 1 3
0 2
0
0 0 53360 0
0
5 GND17
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3524 0 0
2
44519.9 44
0
6 1K RAM
79 1672 404 0 20 41
0 2 2 2 2 2 2 2 67 66
65 117 118 119 120 75 76 77 87 52
10
0
0 0 4848 0
5 RAM1K
-17 -19 18 -11
3 U12
-11 -70 10 -62
0
16 DVCC=22;DGND=11;
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 512 1 0 0 0
1 U
629 0 0
2
44519.9 45
0
9 Inverter~
13 762 176 0 2 22
0 41 63
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
3691 0 0
2
5.90009e-315 5.51416e-315
0
9 Terminal~
194 86 218 0 1 3
0 30
0
0 0 49520 180
7 output3
-46 4 3 12
3 T60
-10 -32 11 -24
0
8 output3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9520 0 0
2
5.90009e-315 5.51481e-315
0
12 Hex Display~
7 89 179 0 16 19
10 31 32 30 33 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3928 0 0
2
5.90009e-315 5.51545e-315
0
9 Terminal~
194 98 218 0 1 3
0 31
0
0 0 49520 180
7 output1
7 -11 56 -3
3 T57
-10 -32 11 -24
0
8 output1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7668 0 0
2
5.90009e-315 5.5161e-315
0
9 Terminal~
194 92 218 0 1 3
0 32
0
0 0 49520 180
7 output2
3 5 52 13
3 T58
-10 -32 11 -24
0
8 output2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5574 0 0
2
5.90009e-315 5.51675e-315
0
9 Terminal~
194 80 218 0 1 3
0 33
0
0 0 49520 180
7 output4
-56 -9 -7 -1
3 T59
-10 -32 11 -24
0
8 output4;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8529 0 0
2
5.90009e-315 5.5174e-315
0
6 74LS83
105 547 569 0 14 29
0 2 2 39 34 2 21 88 22 2
35 36 38 37 121
0
0 0 4848 0
6 74LS83
-21 -60 21 -52
2 U4
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3991 0 0
2
5.90009e-315 5.51804e-315
0
9 Inverter~
13 420 587 0 2 22
0 20 88
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
4208 0 0
2
5.90009e-315 5.51869e-315
0
9 Terminal~
194 489 580 0 1 3
0 21
0
0 0 49520 90
7 clinha1
-55 -7 -6 1
3 T23
-10 -32 11 -24
0
8 clinha1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3445 0 0
2
5.90009e-315 5.51934e-315
0
9 Terminal~
194 393 589 0 1 3
0 20
0
0 0 49520 90
7 clinha3
-55 -7 -6 1
3 T24
-10 -32 11 -24
0
8 clinha3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8822 0 0
2
5.90009e-315 5.51999e-315
0
9 Terminal~
194 489 598 0 1 3
0 22
0
0 0 49520 90
7 clinha2
-55 -7 -6 1
3 T25
-10 -32 11 -24
0
8 clinha2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
530 0 0
2
5.90009e-315 5.52063e-315
0
7 Ground~
168 506 635 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5715 0 0
2
5.90009e-315 5.52128e-315
0
9 Terminal~
194 483 562 0 1 3
0 34
0
0 0 49520 90
6 clock2
-48 -6 -6 2
3 T26
-10 -32 11 -24
0
7 clock2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7530 0 0
2
5.90009e-315 5.52193e-315
0
9 Terminal~
194 616 561 0 1 3
0 35
0
0 0 49520 270
3 sn3
12 -4 33 4
3 T30
-10 -32 11 -24
0
4 sn3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4777 0 0
2
5.90009e-315 5.52258e-315
0
9 Terminal~
194 616 570 0 1 3
0 36
0
0 0 49520 270
3 sn2
12 -4 33 4
3 T31
-10 -32 11 -24
0
4 sn2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3281 0 0
2
5.90009e-315 5.52322e-315
0
9 Terminal~
194 616 588 0 1 3
0 37
0
0 0 49520 270
3 sn0
12 -4 33 4
3 T32
-10 -32 11 -24
0
4 sn0;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5561 0 0
2
5.90009e-315 5.52387e-315
0
9 Terminal~
194 616 579 0 1 3
0 38
0
0 0 49520 270
3 sn1
12 -4 33 4
3 T33
-10 -32 11 -24
0
4 sn1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9298 0 0
2
5.90009e-315 5.52452e-315
0
9 Terminal~
194 483 553 0 1 3
0 39
0
0 0 49520 90
6 clock3
-48 -6 -6 2
3 T27
-10 -32 11 -24
0
7 clock3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9655 0 0
2
5.90009e-315 5.52517e-315
0
9 Terminal~
194 483 723 0 1 3
0 34
0
0 0 49520 90
6 clock2
-48 -6 -6 2
3 T38
-10 -32 11 -24
0
7 clock2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3170 0 0
2
5.90009e-315 5.52581e-315
0
9 Inverter~
13 516 721 0 2 22
0 34 40
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
36 0 0
2
5.90009e-315 5.52646e-315
0
9 Terminal~
194 584 713 0 1 3
0 40
0
0 0 49520 270
3 se3
12 -4 33 4
3 T37
-10 -32 11 -24
0
4 se3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3767 0 0
2
5.90009e-315 5.52711e-315
0
9 Terminal~
194 584 722 0 1 3
0 40
0
0 0 49520 270
3 se2
12 -4 33 4
3 T36
-10 -32 11 -24
0
4 se2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7237 0 0
2
5.90009e-315 5.52776e-315
0
9 Terminal~
194 584 740 0 1 3
0 39
0
0 0 49520 270
3 se0
12 -4 33 4
3 T35
-10 -32 11 -24
0
4 se0;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
863 0 0
2
5.90009e-315 5.52841e-315
0
9 Terminal~
194 584 731 0 1 3
0 40
0
0 0 49520 270
3 se1
12 -4 33 4
3 T34
-10 -32 11 -24
0
4 se1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3881 0 0
2
5.90009e-315 5.52905e-315
0
9 Terminal~
194 535 741 0 1 3
0 39
0
0 0 49520 90
6 clock3
-48 -6 -6 2
3 T29
-10 -32 11 -24
0
7 clock3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9317 0 0
2
5.90009e-315 5.5297e-315
0
9 Terminal~
194 166 466 0 1 3
0 16
0
0 0 49520 270
5 clock
5 -4 40 4
3 T28
-10 -32 11 -24
0
6 clock;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6556 0 0
2
5.90009e-315 5.53035e-315
0
9 2-In AND~
219 105 549 0 3 22
0 16 41 89
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3726 0 0
2
5.90009e-315 5.531e-315
0
9 Terminal~
194 58 560 0 1 3
0 41
0
0 0 49520 90
5 block
-18 -15 17 -7
3 T62
-10 -32 11 -24
0
6 block;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8183 0 0
2
5.90009e-315 5.53164e-315
0
9 Terminal~
194 777 136 0 1 3
0 41
0
0 0 49520 270
5 block
-31 -19 4 -11
3 T61
-10 -32 11 -24
0
6 block;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7993 0 0
2
5.90009e-315 5.53229e-315
0
5 4013~
219 974 747 0 6 22
0 2 90 25 2 122 31
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U8B
24 -54 45 -46
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 3 0
1 U
7733 0 0
2
5.90009e-315 5.53294e-315
0
7 Ground~
168 1026 760 0 1 3
0 2
0
0 0 53360 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3294 0 0
2
5.90009e-315 5.53359e-315
0
9 Terminal~
194 1067 712 0 1 3
0 31
0
0 0 49520 270
7 output1
3 -7 52 1
3 T56
-10 -32 11 -24
0
8 output1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8743 0 0
2
5.90009e-315 5.53423e-315
0
9 Terminal~
194 938 731 0 1 3
0 25
0
0 0 49520 90
3 set
-35 -6 -14 2
3 T55
-10 -32 11 -24
0
4 set;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3127 0 0
2
5.90009e-315 5.53488e-315
0
5 4013~
219 971 630 0 6 22
0 2 91 25 2 123 32
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U8A
24 -54 45 -46
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 3 0
1 U
3312 0 0
2
5.90009e-315 5.53553e-315
0
7 Ground~
168 1023 643 0 1 3
0 2
0
0 0 53360 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6715 0 0
2
5.90009e-315 5.53618e-315
0
9 Terminal~
194 1064 595 0 1 3
0 32
0
0 0 49520 270
7 output2
3 -7 52 1
3 T54
-10 -32 11 -24
0
8 output2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
523 0 0
2
5.90009e-315 5.53682e-315
0
9 Terminal~
194 921 614 0 1 3
0 25
0
0 0 49520 90
3 set
-35 -6 -14 2
3 T53
-10 -32 11 -24
0
4 set;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3831 0 0
2
5.90009e-315 5.53747e-315
0
5 4013~
219 968 519 0 6 22
0 2 92 25 2 124 30
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U7B
24 -54 45 -46
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 2 0
1 U
7292 0 0
2
5.90009e-315 5.53812e-315
0
7 Ground~
168 1020 532 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6123 0 0
2
5.90009e-315 5.53877e-315
0
9 Terminal~
194 1061 484 0 1 3
0 30
0
0 0 49520 270
7 output3
3 -7 52 1
3 T52
-10 -32 11 -24
0
8 output3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3194 0 0
2
5.90009e-315 5.53941e-315
0
9 Terminal~
194 920 503 0 1 3
0 25
0
0 0 49520 90
3 set
-35 -6 -14 2
3 T49
-10 -32 11 -24
0
4 set;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4222 0 0
2
5.90009e-315 5.54006e-315
0
9 Terminal~
194 912 390 0 1 3
0 25
0
0 0 49520 90
3 set
-35 -6 -14 2
3 T51
-10 -32 11 -24
0
4 set;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8263 0 0
2
5.90009e-315 5.54071e-315
0
9 Terminal~
194 1059 371 0 1 3
0 33
0
0 0 49520 270
7 output4
3 -7 52 1
3 T48
-10 -32 11 -24
0
8 output4;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7890 0 0
2
5.90009e-315 5.54136e-315
0
7 Ground~
168 1018 419 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7723 0 0
2
5.90009e-315 5.542e-315
0
5 4013~
219 966 406 0 6 22
0 2 93 25 2 125 33
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U7A
24 -54 45 -46
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 2 0
1 U
8516 0 0
2
5.90009e-315 5.54265e-315
0
9 Terminal~
194 741 544 0 1 3
0 42
0
0 0 49520 90
6 linha4
-47 -15 -5 -7
3 T47
-10 -32 11 -24
0
7 linha4;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3440 0 0
2
5.90009e-315 5.5433e-315
0
9 Terminal~
194 741 616 0 1 3
0 39
0
0 0 49520 90
3 se0
-34 -6 -13 2
3 T46
-10 -32 11 -24
0
4 se0;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5588 0 0
2
5.90009e-315 5.54395e-315
0
9 Terminal~
194 741 607 0 1 3
0 37
0
0 0 49520 90
3 sn0
-34 -6 -13 2
3 T45
-10 -32 11 -24
0
4 sn0;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5857 0 0
2
5.90009e-315 5.54459e-315
0
9 Terminal~
194 741 598 0 1 3
0 40
0
0 0 49520 90
3 se1
-35 -6 -14 2
3 T44
-10 -32 11 -24
0
4 se1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
755 0 0
2
5.90009e-315 5.54524e-315
0
9 Terminal~
194 741 589 0 1 3
0 38
0
0 0 49520 90
3 sn1
-35 -6 -14 2
3 T43
-10 -32 11 -24
0
4 sn1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3400 0 0
2
5.90009e-315 5.54589e-315
0
9 Terminal~
194 741 580 0 1 3
0 40
0
0 0 49520 90
3 se2
-36 -5 -15 3
3 T42
-10 -32 11 -24
0
4 se2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9446 0 0
2
5.90009e-315 5.54654e-315
0
9 Terminal~
194 741 571 0 1 3
0 36
0
0 0 49520 90
3 sn2
-35 -6 -14 2
3 T41
-10 -32 11 -24
0
4 sn2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5210 0 0
2
5.90009e-315 5.54719e-315
0
9 Terminal~
194 741 562 0 1 3
0 40
0
0 0 49520 90
3 se3
-36 -6 -15 2
3 T40
-10 -32 11 -24
0
4 se3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8400 0 0
2
5.90009e-315 5.54783e-315
0
9 Terminal~
194 741 553 0 1 3
0 35
0
0 0 49520 90
3 sn3
-35 -6 -14 2
3 T39
-10 -32 11 -24
0
4 sn3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5909 0 0
2
5.90009e-315 5.54848e-315
0
7 Ground~
168 739 645 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7312 0 0
2
5.90009e-315 5.54913e-315
0
7 74LS157
122 784 578 0 14 29
0 42 35 40 36 40 38 40 37 39
2 93 92 91 90
0
0 0 4848 0
7 74LS157
-24 -60 25 -52
2 U6
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
3838 0 0
2
5.90009e-315 5.54978e-315
0
7 Ground~
168 711 201 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6348 0 0
2
5.90009e-315 5.55042e-315
0
9 Terminal~
194 600 196 0 1 3
0 39
0
0 0 49520 90
6 clock3
-50 -5 -8 3
3 T22
-10 -32 11 -24
0
7 clock3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3466 0 0
2
5.90009e-315 5.55107e-315
0
9 Terminal~
194 600 205 0 1 3
0 34
0
0 0 49520 90
6 clock2
-49 -5 -7 3
3 T21
-10 -32 11 -24
0
7 clock2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3713 0 0
2
5.90009e-315 5.55172e-315
0
9 Terminal~
194 600 169 0 1 3
0 43
0
0 0 49520 90
7 coluna3
-55 -7 -6 1
3 T20
-10 -32 11 -24
0
8 coluna3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4635 0 0
2
5.90009e-315 5.55237e-315
0
9 Terminal~
194 600 178 0 1 3
0 44
0
0 0 49520 90
7 coluna2
-55 -7 -6 1
3 T19
-10 -32 11 -24
0
8 coluna2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4444 0 0
2
5.90009e-315 5.55301e-315
0
9 Terminal~
194 600 187 0 1 3
0 45
0
0 0 49520 90
7 coluna1
-55 -7 -6 1
3 T18
-10 -32 11 -24
0
8 coluna1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3328 0 0
2
5.90009e-315 5.55366e-315
0
9 Terminal~
194 514 366 0 1 3
0 43
0
0 0 49520 180
7 coluna3
4 -7 53 1
3 T17
-10 -32 11 -24
0
8 coluna3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
312 0 0
2
5.90009e-315 5.55398e-315
0
9 Terminal~
194 433 368 0 1 3
0 44
0
0 0 49520 180
7 coluna2
4 -7 53 1
3 T16
-10 -32 11 -24
0
8 coluna2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8412 0 0
2
5.90009e-315 5.55431e-315
0
9 Terminal~
194 343 403 0 1 3
0 45
0
0 0 49520 180
7 coluna1
4 -7 53 1
3 T15
-10 -32 11 -24
0
8 coluna1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6185 0 0
2
5.90009e-315 5.55463e-315
0
7 74LS153
119 665 194 0 14 29
0 64 43 44 45 39 34 126 127 128
129 2 130 41 131
0
0 0 4848 0
7 74LS153
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 512 1 0 0 0
1 U
6455 0 0
2
5.90009e-315 5.55496e-315
0
9 Terminal~
194 282 532 0 1 3
0 39
0
0 0 49520 270
6 clock3
2 -4 44 4
3 T14
-10 -32 11 -24
0
7 clock3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3265 0 0
2
5.90009e-315 5.55528e-315
0
9 Terminal~
194 282 541 0 1 3
0 34
0
0 0 49520 270
6 clock2
2 -5 44 3
3 T13
-10 -32 11 -24
0
7 clock2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9479 0 0
2
5.90009e-315 5.5556e-315
0
2 +V
167 343 55 0 1 3
0 94
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9330 0 0
2
5.90009e-315 5.55593e-315
0
9 Terminal~
194 206 155 0 1 3
0 46
0
0 0 49520 90
6 linha1
-12 -17 30 -9
3 T12
-10 -32 11 -24
0
7 linha1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6531 0 0
2
5.90009e-315 5.55625e-315
0
9 Terminal~
194 206 218 0 1 3
0 47
0
0 0 49520 90
6 linha2
-21 -15 21 -7
3 T11
-10 -32 11 -24
0
7 linha2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9789 0 0
2
5.90009e-315 5.55657e-315
0
9 Terminal~
194 204 281 0 1 3
0 48
0
0 0 49520 90
6 linha3
-21 -15 21 -7
3 T10
-10 -32 11 -24
0
7 linha3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8535 0 0
2
5.90009e-315 5.5569e-315
0
9 Terminal~
194 205 344 0 1 3
0 42
0
0 0 49520 90
6 linha4
-21 -15 21 -7
2 T9
-7 -32 7 -24
0
7 linha4;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3512 0 0
2
5.90009e-315 5.55722e-315
0
9 Terminal~
194 233 646 0 1 3
0 47
0
0 0 49520 270
6 linha2
2 -5 44 3
2 T8
-7 -32 7 -24
0
7 linha2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9912 0 0
2
5.90009e-315 5.55755e-315
0
9 Terminal~
194 233 655 0 1 3
0 46
0
0 0 49520 270
6 linha1
2 -4 44 4
2 T7
-7 -32 7 -24
0
7 linha1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3212 0 0
2
5.90009e-315 5.55787e-315
0
9 Terminal~
194 233 637 0 1 3
0 48
0
0 0 49520 270
6 linha3
2 -4 44 4
2 T6
-7 -32 7 -24
0
7 linha3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8247 0 0
2
5.90009e-315 5.55819e-315
0
9 Terminal~
194 233 628 0 1 3
0 42
0
0 0 49520 270
6 linha4
2 -4 44 4
2 T5
-7 -32 7 -24
0
7 linha4;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3947 0 0
2
5.90009e-315 5.55852e-315
0
9 Terminal~
194 98 647 0 1 3
0 24
0
0 0 49520 90
6 clock0
-48 -4 -6 4
2 T4
-7 -32 7 -24
0
7 clock0;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4251 0 0
2
5.90009e-315 5.55884e-315
0
9 Terminal~
194 98 638 0 1 3
0 23
0
0 0 49520 90
6 clock1
-45 -6 -3 2
2 T3
-7 -32 7 -24
0
7 clock1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
938 0 0
2
5.90009e-315 5.55917e-315
0
9 Terminal~
194 282 559 0 1 3
0 24
0
0 0 49520 270
6 clock0
2 -5 44 3
2 T2
-7 -32 7 -24
0
7 clock0;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3536 0 0
2
5.90009e-315 5.55949e-315
0
9 Terminal~
194 282 550 0 1 3
0 23
0
0 0 49520 270
6 clock1
2 -4 44 4
2 T1
-7 -32 7 -24
0
7 clock1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7643 0 0
2
5.90009e-315 5.55981e-315
0
7 Ground~
168 135 721 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3236 0 0
2
5.90009e-315 5.56014e-315
0
7 Pulser~
4 74 474 0 10 12
0 132 133 16 18 0 0 10 10 7
8
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3903 0 0
2
5.90009e-315 5.56046e-315
0
14 NO PushButton~
191 477 317 0 2 5
0 43 42
0
0 0 4208 0
0
3 S15
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3968 0 0
2
5.90009e-315 5.56078e-315
0
14 NO PushButton~
191 396 316 0 2 5
0 44 42
0
0 0 4208 0
0
3 S14
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3106 0 0
2
5.90009e-315 5.56111e-315
0
14 NO PushButton~
191 314 316 0 2 5
0 45 42
0
0 0 4208 0
0
3 S13
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3223 0 0
2
5.90009e-315 5.56143e-315
0
14 NO PushButton~
191 478 254 0 2 5
0 43 48
0
0 0 4208 0
0
3 S11
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
6341 0 0
2
5.90009e-315 5.56176e-315
0
14 NO PushButton~
191 397 253 0 2 5
0 44 48
0
0 0 4208 0
0
3 S10
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
4627 0 0
2
5.90009e-315 5.56208e-315
0
14 NO PushButton~
191 315 253 0 2 5
0 45 48
0
0 0 4208 0
0
2 S9
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
6952 0 0
2
5.90009e-315 5.5624e-315
0
14 NO PushButton~
191 478 191 0 2 5
0 43 47
0
0 0 4208 0
0
2 S7
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3974 0 0
2
5.90009e-315 5.56273e-315
0
14 NO PushButton~
191 397 190 0 2 5
0 44 47
0
0 0 4208 0
0
2 S5
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
4630 0 0
2
5.90009e-315 5.56305e-315
0
14 NO PushButton~
191 315 190 0 2 5
0 45 47
0
0 0 4208 0
0
2 S4
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
5705 0 0
2
5.90009e-315 5.56337e-315
0
14 NO PushButton~
191 477 128 0 2 5
0 43 46
0
0 0 4208 0
0
2 S3
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
8423 0 0
2
5.90009e-315 5.5637e-315
0
14 NO PushButton~
191 396 127 0 2 5
0 44 46
0
0 0 4208 0
0
2 S2
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
6486 0 0
2
5.90009e-315 5.56402e-315
0
14 NO PushButton~
191 314 127 0 2 5
0 45 46
0
0 0 4208 0
0
2 S1
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3367 0 0
2
5.90009e-315 5.56435e-315
0
9 Resistor~
219 433 90 0 4 5
0 44 94 0 1
0
0 0 880 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7389 0 0
2
5.90009e-315 5.56467e-315
0
9 Resistor~
219 514 89 0 4 5
0 43 94 0 1
0
0 0 880 90
2 1k
8 0 22 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6782 0 0
2
5.90009e-315 5.56499e-315
0
9 Resistor~
219 343 89 0 4 5
0 45 94 0 1
0
0 0 880 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5728 0 0
2
5.90009e-315 5.56532e-315
0
272
1 1 2 0 0 12288 0 99 9 0 0 4
1710 1238
1710 1224
1679 1224
1679 1315
2 1 49 0 0 4224 0 99 10 0 0 3
1686 1259
1663 1259
1663 1244
1 4 3 0 0 4096 0 11 99 0 0 2
1710 1313
1710 1301
1 1 28 0 0 8192 0 101 12 0 0 3
1792 1258
1792 1262
1843 1262
1 1 4 0 0 8192 0 1 13 0 0 3
1948 1350
1948 1352
1973 1352
1 2 50 0 0 4224 0 14 114 0 0 3
1293 955
1293 1007
1342 1007
1 1 5 0 0 4096 0 57 15 0 0 2
1130 1625
1177 1625
1 3 17 0 0 4096 0 52 54 0 0 2
1220 1673
1168 1673
1 0 2 0 0 0 0 16 0 0 16 3
1603 997
1592 997
1592 1033
3 1 51 0 0 8320 0 16 2 0 0 4
1603 1015
1586 1015
1586 965
1572 965
1 2 5 0 0 0 0 23 16 0 0 2
1578 1006
1609 1006
1 4 10 0 0 4096 0 22 16 0 0 2
1578 1024
1609 1024
8 0 2 0 0 0 0 16 0 0 16 2
1609 1060
1592 1060
7 0 2 0 0 0 0 16 0 0 16 2
1609 1051
1592 1051
6 0 2 0 0 0 0 16 0 0 16 2
1609 1042
1592 1042
5 1 2 0 0 0 0 16 21 0 0 3
1609 1033
1592 1033
1592 1111
1 12 6 0 0 4096 0 17 16 0 0 2
1687 1042
1673 1042
1 11 9 0 0 4224 0 20 16 0 0 2
1739 1033
1673 1033
1 14 8 0 0 4096 0 19 16 0 0 2
1687 1060
1673 1060
1 13 7 0 0 4096 0 18 16 0 0 2
1687 1051
1673 1051
2 19 52 0 0 8320 0 24 136 0 0 4
1690 297
1724 297
1724 368
1710 368
1 3 6 0 0 4224 0 27 26 0 0 2
1684 746
1684 721
1 2 7 0 0 0 0 28 26 0 0 2
1690 733
1690 721
1 1 8 0 0 0 0 29 26 0 0 2
1696 721
1696 721
1 3 13 0 0 4096 0 32 33 0 0 2
1600 748
1600 723
1 2 12 0 0 4096 0 31 33 0 0 2
1606 735
1606 723
1 1 11 0 0 0 0 30 33 0 0 2
1612 723
1612 723
1 0 10 0 0 0 0 34 0 0 161 2
1762 154
1741 154
1 -208000 53 0 0 8320 0 35 0 0 128 3
2154 368
2154 430
2062 430
2 -207999 54 0 0 8320 0 35 0 0 128 3
2148 368
2148 416
2062 416
-207998 3 55 0 0 4224 0 0 35 128 0 3
2062 403
2142 403
2142 368
4 -207997 56 0 0 8320 0 35 0 0 128 3
2136 368
2136 391
2062 391
2 4 57 0 0 8320 0 45 39 0 0 4
1713 1532
1702 1532
1702 1554
1697 1554
3 1 8 0 0 4224 0 39 38 0 0 2
1651 1563
1634 1563
2 1 7 0 0 4224 0 39 37 0 0 2
1652 1554
1634 1554
1 1 6 0 0 0 0 39 36 0 0 2
1651 1545
1634 1545
1 3 15 0 0 4224 0 44 45 0 0 2
1796 1523
1758 1523
1 1 16 0 0 4096 0 45 46 0 0 2
1713 1514
1690 1514
1 3 3 0 0 4224 0 43 41 0 0 2
1795 1467
1757 1467
1 2 14 0 0 4096 0 42 41 0 0 2
1690 1476
1712 1476
1 1 10 0 0 0 0 41 40 0 0 2
1712 1458
1689 1458
6 3 58 0 0 4224 0 87 50 0 0 3
1491 557
1276 557
1276 604
1 0 59 0 0 4096 0 50 0 0 83 2
1267 649
1267 656
1 1 6 0 0 128 0 48 49 0 0 2
1276 730
1276 711
1 2 9 0 0 128 0 47 49 0 0 2
1294 731
1294 711
2 3 60 0 0 4224 0 50 49 0 0 2
1285 649
1285 665
2 3 61 0 0 4224 0 51 114 0 0 4
1396 962
1311 962
1311 1016
1336 1016
11 1 62 0 0 8320 0 114 51 0 0 4
1406 1034
1446 1034
1446 962
1432 962
1 2 10 0 0 4224 0 53 54 0 0 2
1047 1682
1123 1682
0 1 5 0 0 0 0 0 54 52 0 3
1110 1625
1110 1664
1123 1664
1 1 14 0 0 0 0 55 56 0 0 2
1045 1616
1061 1616
3 1 5 0 0 0 0 56 57 0 0 2
1106 1625
1130 1625
1 2 18 0 0 4096 0 58 56 0 0 2
1045 1634
1061 1634
14 1 21 0 0 4096 0 68 61 0 0 2
219 690
221 690
13 1 22 0 0 4096 0 68 62 0 0 2
219 681
221 681
12 1 20 0 0 4224 0 68 60 0 0 2
219 672
221 672
11 1 19 0 0 4224 0 68 59 0 0 2
219 663
221 663
6 0 2 0 0 0 0 68 0 0 267 2
143 690
135 690
1 5 24 0 0 4096 0 64 68 0 0 2
107 681
149 681
1 4 23 0 0 4096 0 63 68 0 0 2
107 672
149 672
1 2 16 0 0 4096 0 65 66 0 0 2
784 193
809 193
3 1 25 0 0 4224 0 66 70 0 0 2
854 184
906 184
2 1 63 0 0 8320 0 137 66 0 0 3
783 176
783 175
809 175
1 1 64 0 0 8320 0 202 67 0 0 3
633 158
617 158
617 136
10 1 46 0 0 4096 0 68 211 0 0 2
219 654
221 654
9 1 47 0 0 4096 0 68 210 0 0 2
219 645
221 645
8 1 48 0 0 4096 0 68 212 0 0 2
219 636
221 636
7 1 42 0 0 4096 0 68 213 0 0 2
219 627
221 627
10 -1535 65 0 0 4224 0 136 0 0 75 2
1640 449
1596 449
9 -1534 66 0 0 4224 0 136 0 0 75 2
1640 440
1596 440
8 -1533 67 0 0 4224 0 136 0 0 75 2
1640 431
1596 431
13 -1535 65 0 0 0 0 87 0 0 75 2
1555 566
1596 566
12 -1534 66 0 0 0 0 87 0 0 75 2
1555 557
1596 557
11 -1533 67 0 0 0 0 87 0 0 75 2
1555 548
1596 548
-95129 0 1 0 0 4128 0 0 0 0 0 2
1596 352
1596 624
0 1 59 0 0 4224 0 0 77 83 0 3
1331 656
1403 656
1403 651
1 2 9 0 0 0 0 80 78 0 0 2
1430 728
1430 712
1 1 8 0 0 128 0 79 78 0 0 2
1412 728
1412 712
2 3 68 0 0 4224 0 77 78 0 0 2
1421 651
1421 666
1 2 9 0 0 0 0 76 72 0 0 2
1358 726
1358 710
1 1 7 0 0 128 0 75 72 0 0 2
1340 726
1340 710
1 1 10 0 0 128 0 71 74 0 0 2
1175 656
1206 656
2 1 59 0 0 4224 0 74 73 0 0 3
1242 656
1331 656
1331 649
2 3 69 0 0 4224 0 73 72 0 0 2
1349 649
1349 664
3 7 70 0 0 8320 0 73 87 0 0 3
1340 604
1340 566
1491 566
7 0 2 0 0 0 0 136 0 0 167 2
1640 422
1624 422
1 14 11 0 0 4096 0 83 114 0 0 2
1419 1061
1406 1061
1 13 12 0 0 4096 0 82 114 0 0 2
1419 1052
1406 1052
1 12 13 0 0 0 0 81 114 0 0 2
1419 1043
1406 1043
14 0 2 0 0 0 0 87 0 0 97 4
1555 593
1565 593
1565 611
1475 611
1 2 13 0 0 4224 0 84 87 0 0 2
1458 521
1491 521
1 3 12 0 0 4224 0 85 87 0 0 2
1458 530
1491 530
1 4 11 0 0 4224 0 86 87 0 0 2
1458 539
1491 539
3 8 71 0 0 8320 0 77 87 0 0 3
1412 606
1412 575
1491 575
9 0 2 0 0 0 0 87 0 0 97 2
1491 593
1475 593
5 0 2 0 0 0 0 87 0 0 97 2
1491 548
1475 548
1 1 2 0 0 8320 0 87 88 0 0 3
1491 512
1475 512
1475 658
4 1 18 0 0 4096 0 219 91 0 0 4
104 474
129 474
129 485
154 485
2 2 72 0 0 4224 0 92 90 0 0 2
1347 1504
1363 1504
3 1 26 0 0 4096 0 90 93 0 0 2
1408 1495
1452 1495
1 1 9 0 0 0 0 94 92 0 0 3
1267 1502
1267 1504
1311 1504
1 1 18 0 0 4224 0 90 95 0 0 2
1363 1486
1304 1486
3 1 27 0 0 4096 0 89 98 0 0 2
1103 1495
1134 1495
1 2 9 0 0 0 0 97 89 0 0 3
1035 1503
1035 1504
1058 1504
1 1 16 0 0 4224 0 89 96 0 0 2
1058 1486
1000 1486
6 1 28 0 0 4224 0 99 101 0 0 3
1734 1259
1792 1259
1792 1258
3 1 15 0 0 4224 0 99 100 0 0 3
1686 1277
1644 1277
1644 1276
1 1 2 0 0 0 0 102 107 0 0 4
1400 1238
1400 1220
1371 1220
1371 1331
6 1 29 0 0 4224 0 102 106 0 0 3
1424 1259
1482 1259
1482 1258
1 4 26 0 0 4224 0 105 102 0 0 3
1332 1313
1400 1313
1400 1301
3 1 27 0 0 4224 0 102 104 0 0 3
1376 1277
1299 1277
1299 1275
1 2 73 0 0 8320 0 103 102 0 0 3
1339 1256
1339 1259
1376 1259
1 1 2 0 0 0 0 113 108 0 0 4
1105 1239
1105 1221
1076 1221
1076 1332
6 1 14 0 0 4224 0 113 109 0 0 3
1129 1260
1187 1260
1187 1259
1 4 5 0 0 4224 0 110 113 0 0 3
1037 1314
1105 1314
1105 1302
3 1 4 0 0 4224 0 113 111 0 0 3
1081 1278
1004 1278
1004 1276
1 2 74 0 0 8320 0 112 113 0 0 3
1044 1257
1044 1260
1081 1260
1 1 17 0 0 4224 0 114 116 0 0 2
1342 998
1260 998
0 4 2 0 0 0 0 0 114 123 0 3
1326 1034
1326 1025
1342 1025
8 0 2 0 0 0 0 114 0 0 123 2
1342 1061
1325 1061
7 0 2 0 0 0 0 114 0 0 123 2
1342 1052
1325 1052
6 0 2 0 0 0 0 114 0 0 123 2
1342 1043
1325 1043
5 1 2 0 0 0 0 114 115 0 0 3
1342 1034
1325 1034
1325 1107
13 -207997 56 0 0 128 0 134 0 0 128 2
1991 321
2062 321
14 -207998 55 0 0 128 0 134 0 0 128 2
1991 330
2062 330
15 -207999 54 0 0 128 0 134 0 0 128 2
1991 339
2062 339
16 -208000 53 0 0 128 0 134 0 0 128 2
1991 348
2062 348
-13308169 0 1 0 0 4256 0 0 0 0 0 2
2062 138
2062 707
1 1 4 0 0 128 0 25 24 0 0 2
1619 297
1654 297
18 0 10 0 0 12416 0 134 0 0 161 4
1991 276
2002 276
2002 217
1741 217
1 17 2 0 0 0 0 117 134 0 0 3
1904 296
1904 276
1921 276
5 -3261 75 0 0 4096 0 134 0 0 160 2
1927 321
1823 321
6 -3262 76 0 0 4096 0 134 0 0 160 2
1927 330
1823 330
7 -3263 77 0 0 4096 0 134 0 0 160 2
1927 339
1823 339
3 0 78 0 0 4096 0 118 0 0 138 2
2517 207
2435 207
3 0 78 0 0 0 0 125 0 0 138 2
2514 349
2435 349
3 0 78 0 0 0 0 129 0 0 138 2
2514 497
2435 497
1 3 78 0 0 8320 0 7 133 0 0 4
2422 149
2435 149
2435 637
2517 637
6 1 79 0 0 4224 0 133 130 0 0 2
2565 619
2611 619
4 1 2 0 0 0 0 133 131 0 0 2
2541 661
2541 673
1 1 2 0 0 0 0 133 132 0 0 4
2541 598
2541 559
2641 559
2641 572
1 2 80 0 0 4224 0 6 133 0 0 2
2487 619
2517 619
6 1 81 0 0 4224 0 129 126 0 0 2
2562 479
2608 479
4 1 2 0 0 0 0 129 127 0 0 2
2538 521
2538 533
1 1 2 0 0 0 0 129 128 0 0 4
2538 458
2538 419
2645 419
2645 428
1 2 82 0 0 4224 0 5 129 0 0 2
2484 479
2514 479
6 1 83 0 0 4224 0 125 122 0 0 2
2562 331
2610 331
4 1 2 0 0 0 0 125 123 0 0 2
2538 373
2538 387
1 1 2 0 0 0 0 125 124 0 0 4
2538 310
2538 273
2645 273
2645 284
1 2 84 0 0 4224 0 4 125 0 0 2
2482 331
2514 331
6 1 85 0 0 4224 0 118 121 0 0 2
2565 189
2611 189
4 1 2 0 0 0 0 118 120 0 0 2
2541 231
2541 243
1 1 2 0 0 0 0 118 119 0 0 4
2541 168
2541 129
2647 129
2647 143
1 2 86 0 0 4224 0 3 118 0 0 2
2487 189
2517 189
8 -3264 87 0 0 4096 0 134 0 0 160 2
1927 348
1823 348
15 -3261 75 0 0 4224 0 136 0 0 160 2
1704 422
1823 422
16 -3262 76 0 0 4224 0 136 0 0 160 2
1704 431
1823 431
17 -3263 77 0 0 4224 0 136 0 0 160 2
1704 440
1823 440
18 -3264 87 0 0 4224 0 136 0 0 160 2
1704 449
1823 449
-846037834 0 1 0 0 32 0 0 0 0 0 2
1823 140
1823 709
1 20 10 0 0 0 0 8 136 0 0 4
1608 154
1741 154
1741 377
1710 377
6 0 2 0 0 0 0 136 0 0 167 2
1640 413
1624 413
5 0 2 0 0 0 0 136 0 0 167 2
1640 404
1624 404
4 0 2 0 0 0 0 136 0 0 167 2
1640 395
1624 395
3 0 2 0 0 0 0 136 0 0 167 2
1640 386
1624 386
2 0 2 0 0 0 0 136 0 0 167 2
1640 377
1624 377
1 1 2 0 0 0 0 136 135 0 0 3
1640 368
1624 368
1624 473
0 1 40 0 0 8192 0 0 160 189 0 3
555 721
555 730
572 730
1 3 30 0 0 0 0 138 139 0 0 2
86 203
86 203
1 4 33 0 0 0 0 142 139 0 0 2
80 203
80 203
1 2 32 0 0 0 0 141 139 0 0 2
92 203
92 203
1 1 31 0 0 0 0 140 139 0 0 2
98 203
98 203
2 0 2 0 0 0 0 143 0 0 180 2
515 542
506 542
4 1 34 0 0 4096 0 143 149 0 0 2
515 560
494 560
1 3 39 0 0 4096 0 154 143 0 0 2
494 551
515 551
1 13 37 0 0 4224 0 152 143 0 0 2
604 587
579 587
1 12 38 0 0 4224 0 153 143 0 0 2
604 578
579 578
1 11 36 0 0 4224 0 151 143 0 0 2
604 569
579 569
1 10 35 0 0 4224 0 150 143 0 0 2
604 560
579 560
1 0 2 0 0 0 0 143 0 0 182 3
515 533
506 533
506 569
9 0 2 0 0 0 0 143 0 0 182 2
515 614
506 614
5 1 2 0 0 0 0 143 148 0 0 3
515 569
506 569
506 629
1 8 22 0 0 4224 0 147 143 0 0 2
500 596
515 596
2 7 88 0 0 4224 0 144 143 0 0 2
441 587
515 587
1 1 20 0 0 0 0 146 144 0 0 2
404 587
405 587
1 6 21 0 0 4224 0 145 143 0 0 2
500 578
515 578
1 1 34 0 0 0 0 155 156 0 0 2
494 721
501 721
1 1 39 0 0 4096 0 159 161 0 0 2
572 739
546 739
1 2 40 0 0 4224 0 158 156 0 0 2
572 721
537 721
1 0 40 0 0 0 0 157 0 0 189 3
572 712
548 712
548 721
0 1 16 0 0 0 0 0 162 193 0 2
117 465
154 465
3 3 89 0 0 4224 0 163 69 0 0 2
126 549
153 549
1 3 16 0 0 0 0 163 219 0 0 6
81 540
63 540
63 514
117 514
117 465
98 465
1 2 41 0 0 4096 0 164 163 0 0 2
69 558
81 558
0 1 41 0 0 8192 0 0 165 227 0 3
721 176
721 135
765 135
14 2 90 0 0 8320 0 192 166 0 0 4
816 614
873 614
873 711
950 711
13 2 91 0 0 4224 0 192 170 0 0 3
816 596
947 596
947 594
2 12 92 0 0 8320 0 174 192 0 0 4
944 483
873 483
873 578
816 578
11 2 93 0 0 8320 0 192 181 0 0 4
816 560
864 560
864 370
942 370
1 3 25 0 0 0 0 169 166 0 0 2
949 729
950 729
6 1 31 0 0 4224 0 166 168 0 0 2
998 711
1055 711
1 1 2 0 0 0 0 166 167 0 0 3
974 690
1026 690
1026 754
4 1 2 0 0 0 0 166 167 0 0 3
974 753
974 754
1026 754
1 3 25 0 0 0 0 173 170 0 0 2
932 612
947 612
6 1 32 0 0 4224 0 170 172 0 0 2
995 594
1052 594
1 1 2 0 0 0 0 170 171 0 0 3
971 573
1023 573
1023 637
4 1 2 0 0 0 0 170 171 0 0 3
971 636
971 637
1023 637
1 3 25 0 0 0 0 177 174 0 0 2
931 501
944 501
6 1 30 0 0 4224 0 174 176 0 0 2
992 483
1049 483
1 1 2 0 0 0 0 174 175 0 0 3
968 462
1020 462
1020 526
4 1 2 0 0 0 0 174 175 0 0 3
968 525
968 526
1020 526
1 3 25 0 0 0 0 178 181 0 0 2
923 388
942 388
6 1 33 0 0 4224 0 181 179 0 0 2
990 370
1047 370
1 1 2 0 0 0 0 181 180 0 0 3
966 349
1018 349
1018 413
4 1 2 0 0 0 0 181 180 0 0 3
966 412
966 413
1018 413
1 1 42 0 0 0 0 182 192 0 0 2
752 542
752 542
1 8 37 0 0 0 0 184 192 0 0 2
752 605
752 605
1 9 39 0 0 0 0 183 192 0 0 2
752 614
752 614
1 6 38 0 0 0 0 186 192 0 0 4
752 587
753 587
753 587
752 587
1 7 40 0 0 0 0 185 192 0 0 2
752 596
752 596
1 4 36 0 0 0 0 188 192 0 0 2
752 569
752 569
1 5 40 0 0 0 0 187 192 0 0 2
752 578
752 578
1 2 35 0 0 0 0 190 192 0 0 2
752 551
752 551
1 3 40 0 0 0 0 189 192 0 0 2
752 560
752 560
1 10 2 0 0 0 0 191 192 0 0 3
739 639
739 623
746 623
1 11 2 0 0 0 0 193 202 0 0 3
711 195
711 158
703 158
13 1 41 0 0 4224 0 202 137 0 0 2
697 176
747 176
1 5 39 0 0 0 0 194 202 0 0 2
611 194
633 194
1 6 34 0 0 4096 0 195 202 0 0 2
611 203
633 203
1 2 43 0 0 4096 0 196 202 0 0 2
611 167
633 167
1 3 44 0 0 4096 0 197 202 0 0 2
611 176
633 176
1 4 45 0 0 4096 0 198 202 0 0 2
611 185
633 185
6 1 34 0 0 4224 0 69 204 0 0 2
223 540
270 540
5 1 39 0 0 4224 0 69 203 0 0 2
223 531
270 531
2 0 2 0 0 0 0 69 0 0 236 2
159 540
135 540
0 1 2 0 0 0 0 0 69 267 0 3
135 654
135 531
159 531
2 0 46 0 0 4096 0 231 0 0 266 2
297 135
297 153
2 0 46 0 0 0 0 230 0 0 266 2
379 135
379 153
2 0 47 0 0 4096 0 228 0 0 265 2
298 198
298 216
2 0 47 0 0 0 0 227 0 0 265 2
380 198
380 216
2 0 48 0 0 4096 0 225 0 0 264 2
298 261
298 279
2 0 48 0 0 0 0 224 0 0 264 2
380 261
380 279
2 0 42 0 0 4096 0 222 0 0 263 2
297 324
297 342
2 0 42 0 0 0 0 221 0 0 263 2
379 324
379 342
1 0 43 0 0 0 0 220 0 0 259 2
494 325
514 325
1 0 43 0 0 0 0 223 0 0 259 2
495 262
514 262
1 0 43 0 0 0 0 226 0 0 259 2
495 199
514 199
1 0 44 0 0 0 0 221 0 0 260 2
413 324
433 324
1 0 44 0 0 0 0 224 0 0 260 2
414 261
433 261
1 0 44 0 0 0 0 227 0 0 260 2
414 198
433 198
1 0 45 0 0 0 0 222 0 0 261 2
331 324
343 324
1 0 45 0 0 0 0 225 0 0 261 2
332 261
343 261
1 0 45 0 0 0 0 228 0 0 261 2
332 198
343 198
1 0 43 0 0 0 0 229 0 0 259 2
494 136
514 136
1 0 44 0 0 0 0 230 0 0 260 2
413 135
433 135
1 0 45 0 0 0 0 231 0 0 261 2
331 135
343 135
2 2 94 0 0 8192 0 232 233 0 0 3
433 72
433 71
514 71
2 2 94 0 0 4224 0 234 232 0 0 3
343 71
433 71
433 72
1 1 43 0 0 4224 0 233 199 0 0 2
514 107
514 351
1 1 44 0 0 4224 0 232 200 0 0 2
433 108
433 353
1 1 45 0 0 4224 0 234 201 0 0 2
343 107
343 388
2 1 94 0 0 0 0 234 205 0 0 2
343 71
343 64
1 2 42 0 0 4224 0 209 220 0 0 3
216 342
460 342
460 325
1 2 48 0 0 4224 0 208 223 0 0 3
215 279
461 279
461 262
1 2 47 0 0 4224 0 207 226 0 0 3
217 216
461 216
461 199
1 2 46 0 0 4224 0 206 229 0 0 3
217 153
460 153
460 136
3 1 2 0 0 0 0 68 218 0 0 3
143 654
135 654
135 715
1 2 24 0 0 0 0 214 68 0 0 2
109 645
149 645
1 1 23 0 0 0 0 215 68 0 0 2
109 636
149 636
0 1 24 0 0 0 0 0 216 272 0 2
234 558
270 558
7 1 23 0 0 4224 0 69 217 0 0 2
223 549
270 549
8 4 24 0 0 12416 0 69 69 0 0 6
223 558
234 558
234 575
144 575
144 558
153 558
33
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 154
1856 1459 2423 1563
1863 1465 2415 1545
154 IF write_read AND (modo == 1):  // operacao no clockup
   ddown = 1

IF nclock AND (q > 0):  // operacao no clockup (pr�ximo ap�s mudar q)
   ddup = 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
1637 633 1732 657
1644 638 1724 654
10 quantidade
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1570 632 1633 656
1577 638 1625 654
6 inicio
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
1601 1087 1696 1111
1608 1092 1688 1108
10 quantidade
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 103
1254 411 1465 535
1259 415 1459 511
103 ESCRITA (modo=0)
end = inicio + 7 (se q=8)
    = inicio + q (senao)

LEITURA (modo=1)
end = inicio
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 32
1292 1522 1463 1566
1297 1526 1457 1558
32 clock_down AND q!=8:
   or_down
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 24
1016 1521 1139 1565
1021 1525 1133 1557
24 clock AND q=8:
   or_up
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 122
1266 1614 1509 1758
1271 1618 1503 1730
122 IF !clock AND write_read_out:
   write_read = 0
   IF (modo==0):
      q += 1
   ELSE
      q -= 1
      inicio += 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
1101 1322 1196 1346
1108 1327 1188 1343
10 write/read
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 82
2353 60 2736 102
2365 70 2723 100
82 REGISTRADOR (Entradas tempor�rias com chaves s� pra 
mostrar que t� funcionando)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
55 93 120 132
63 100 111 130
14 * -> E
# -> F
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
397 37 540 61
404 42 532 58
16 matriz de botoes
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
295 93 334 117
302 99 326 115
3 (1)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
381 98 412 122
384 100 408 116
3 (2)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
462 99 493 123
465 101 489 117
3 (3)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
300 162 331 186
303 164 327 180
3 (4)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
382 162 413 186
385 164 409 180
3 (5)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
463 163 494 187
466 165 490 181
3 (6)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
300 225 331 249
303 227 327 243
3 (7)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
382 225 413 249
385 227 409 243
3 (8)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
463 226 494 250
466 228 490 244
3 (9)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
381 288 412 312
384 290 408 306
3 (0)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
462 289 493 313
465 291 489 307
3 (#)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
299 288 330 312
302 290 326 306
3 (*)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
147 428 282 452
150 430 278 446
16 divisao do clock
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
454 479 617 503
459 483 611 499
19 aritmetica para 1-9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 24
437 672 640 696
442 676 634 692
24 aritmetica para *, 0 e #
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 51
675 450 838 514
680 454 832 502
51 multiplex para
escolher entre
as duas aritmeticas
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
915 296 998 340
920 300 992 332
20 "memoria"
de 4 bits
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
64 73 119 97
71 78 111 94
5 saida
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1342 1080 1405 1104
1349 1086 1397 1102
6 inicio
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1401 1323 1472 1347
1408 1329 1464 1345
7 overrun
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
1720 1325 1823 1349
1727 1330 1815 1346
11 ddisponivel
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-06 1e-07 1e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
