CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
200 0 30 150 10
176 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.331203 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
277
13 Logic Switch~
5 646 107 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3406 0 0
2
44521.8 0
0
13 Logic Switch~
5 1102 96 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3132 0 0
2
5.90009e-315 0
0
9 Terminal~
194 1156 315 0 1 3
0 2
0
0 0 49520 180
5 qoito
6 -7 41 1
4 T171
-14 -32 14 -24
0
6 qoito;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3842 0 0
2
44521.8 0
0
9 Terminal~
194 822 304 0 1 3
0 3
0
0 0 49520 180
5 ddout
13 -7 48 1
4 T152
-13 -32 15 -24
0
6 ddout;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6183 0 0
2
44521.8 1
0
14 Logic Display~
6 822 271 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3356 0 0
2
44521.8 2
0
9 Terminal~
194 939 305 0 1 3
0 4
0
0 0 49520 180
5 orout
13 -7 48 1
4 T153
-13 -32 15 -24
0
6 orout;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3525 0 0
2
44521.8 3
0
14 Logic Display~
6 939 269 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3800 0 0
2
44521.8 4
0
9 Terminal~
194 708 108 0 1 3
0 5
0
0 0 49520 270
7 letecla
-42 -13 7 -5
4 T151
-13 -32 15 -24
0
8 letecla;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
346 0 0
2
44521.8 5
0
7 Ground~
168 2355 121 0 1 3
0 6
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3169 0 0
2
44521.8 6
0
9 Terminal~
194 2274 197 0 1 3
0 7
0
0 0 49520 90
5 wrout
-43 -6 -8 2
4 T146
-14 -32 14 -24
0
6 wrout;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4826 0 0
2
44521.8 7
0
9 Terminal~
194 1261 1686 0 1 3
0 8
0
0 0 49520 602
6 mododw
-21 -15 21 -7
4 T144
-14 -32 14 -24
0
7 mododw;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3971 0 0
2
44521.8 8
0
9 Terminal~
194 1594 279 0 1 3
0 7
0
0 0 49520 0
5 wrout
-17 -23 18 -15
4 T129
-14 -32 14 -24
0
6 wrout;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3607 0 0
2
44521.8 9
0
9 Inverter~
13 1646 288 0 2 22
0 7 66
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 11 0
1 U
3506 0 0
2
44521.8 10
0
9 Terminal~
194 1632 645 0 1 3
0 9
0
0 0 49520 270
2 e3
-7 -15 7 -7
4 T168
-13 -32 15 -24
0
3 e3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7829 0 0
2
44521.8 11
0
9 Terminal~
194 1626 657 0 1 3
0 10
0
0 0 49520 270
2 e2
-7 -15 7 -7
4 T169
-13 -32 15 -24
0
3 e2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3890 0 0
2
44521.8 12
0
9 Terminal~
194 1620 670 0 1 3
0 11
0
0 0 49520 270
2 e1
-7 -15 7 -7
4 T170
-13 -32 15 -24
0
3 e1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3126 0 0
2
44521.8 13
0
12 Hex Display~
7 1270 237 0 16 19
10 11 10 9 94 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
3935 0 0
2
44521.8 14
0
9 Terminal~
194 1267 301 0 1 3
0 9
0
0 0 49520 180
2 e3
14 -7 28 1
4 T167
-13 -32 15 -24
0
3 e3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9746 0 0
2
44521.8 15
0
9 Terminal~
194 1273 288 0 1 3
0 10
0
0 0 49520 180
2 e2
14 -7 28 1
4 T166
-13 -32 15 -24
0
3 e2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7330 0 0
2
44521.8 16
0
9 Terminal~
194 1279 276 0 1 3
0 11
0
0 0 49520 180
2 e1
14 -7 28 1
4 T164
-13 -32 15 -24
0
3 e1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3972 0 0
2
44521.8 17
0
9 Terminal~
194 1610 1543 0 1 3
0 2
0
0 0 49520 90
5 qoito
-40 -6 -5 2
4 T115
-14 -32 14 -24
0
6 qoito;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7818 0 0
2
44521.8 18
0
9 Terminal~
194 1610 1570 0 1 3
0 12
0
0 0 49520 90
4 qua1
-37 -6 -9 2
4 T120
-14 -32 14 -24
0
5 qua1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3818 0 0
2
44521.8 19
0
9 Terminal~
194 1610 1561 0 1 3
0 13
0
0 0 49520 90
4 qua2
-37 -6 -9 2
4 T119
-14 -32 14 -24
0
5 qua2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8835 0 0
2
44521.8 20
0
9 Terminal~
194 1610 1552 0 1 3
0 14
0
0 0 49520 90
4 qua3
-37 -6 -9 2
4 T118
-14 -32 14 -24
0
5 qua3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7484 0 0
2
44521.8 21
0
8 4-In OR~
219 1656 1554 0 5 22
0 2 14 13 12 36
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U8A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 3 0
1 U
792 0 0
2
44521.8 22
0
9 Terminal~
194 1548 1723 0 1 3
0 15
0
0 0 49520 270
2 pq
-7 -15 7 -7
4 T163
-14 -32 14 -24
0
3 pq;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3826 0 0
2
44521.8 23
0
5 4071~
219 1477 1721 0 3 22
0 67 8 15
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
7958 0 0
2
44521.8 24
0
9 Terminal~
194 1167 1590 0 1 3
0 16
0
0 0 49520 0
6 wrdown
-21 -22 21 -14
4 T114
-14 -32 14 -24
0
7 wrdown;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6736 0 0
2
44521.8 25
0
9 3-In AND~
219 1410 1634 0 4 22
0 16 70 69 67
0
0 0 624 0
6 74LS11
-21 -28 21 -20
4 GNDA
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 0 0
1 U
3755 0 0
2
44521.8 26
0
7 Ground~
168 900 1320 0 1 3
0 6
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
397 0 0
2
44521.8 27
0
9 Terminal~
194 884 1278 0 1 3
0 17
0
0 0 49520 90
5 clock
-18 4 17 12
4 T165
-14 -32 14 -24
0
6 clock;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5190 0 0
2
44521.8 28
0
9 Terminal~
194 782 1269 0 1 3
0 18
0
0 0 49520 90
7 writeup
-24 -15 25 -7
4 T148
-14 -32 14 -24
0
8 writeup;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9188 0 0
2
44521.8 29
0
9 Terminal~
194 781 1251 0 1 3
0 19
0
0 0 49520 90
6 readup
-21 -15 21 -7
3 T73
-11 -32 10 -24
0
7 readup;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3651 0 0
2
44521.8 30
0
8 2-In OR~
219 835 1258 0 3 22
0 19 18 68
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U19D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
3415 0 0
2
44521.8 31
0
5 4013~
219 935 1294 0 6 22
0 6 68 17 6 95 89
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U15B
21 -54 49 -46
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 15 0
1 U
7597 0 0
2
44521.8 32
0
9 Terminal~
194 1546 71 0 1 3
0 18
0
0 0 49520 90
3 set
-11 -15 10 -7
3 T64
-10 -32 11 -24
0
4 set;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
350 0 0
2
5.90009e-315 5.26354e-315
0
9 Inverter~
13 1373 1677 0 2 22
0 4 69
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U3F
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 11 0
1 U
3153 0 0
2
5.90009e-315 5.30499e-315
0
9 Terminal~
194 1376 1726 0 1 3
0 4
0
0 0 49520 180
5 orout
6 -7 41 1
4 T162
-14 -32 14 -24
0
6 orout;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
634 0 0
2
5.90009e-315 5.32571e-315
0
9 Inverter~
13 1344 1634 0 2 22
0 20 70
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 11 0
1 U
8956 0 0
2
5.90009e-315 5.34643e-315
0
9 Terminal~
194 1288 1636 0 1 3
0 20
0
0 0 49520 90
4 modo
-36 -6 -8 2
3 T60
-11 -32 10 -24
0
5 modo;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3342 0 0
2
5.90009e-315 5.3568e-315
0
14 Logic Display~
6 1091 336 0 1 2
10 21
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3549 0 0
2
5.90009e-315 5.36716e-315
0
9 Terminal~
194 1172 355 0 1 3
0 21
0
0 0 49520 270
5 store
3 -5 38 3
3 T59
-10 -32 11 -24
0
6 store;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9177 0 0
2
5.90009e-315 5.37752e-315
0
9 Terminal~
194 2448 144 0 1 3
0 21
0
0 0 49520 270
5 store
3 -5 38 3
3 T58
-10 -32 11 -24
0
6 store;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3387 0 0
2
5.90009e-315 5.38788e-315
0
9 Terminal~
194 1150 86 0 1 3
0 22
0
0 0 49520 0
6 mreset
-22 -22 20 -14
3 T57
-11 -32 10 -24
0
7 mreset;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
351 0 0
2
5.90009e-315 5.39306e-315
0
9 Terminal~
194 1586 920 0 1 3
0 22
0
0 0 49520 0
6 mreset
-22 -22 20 -14
3 T57
-11 -32 10 -24
0
7 mreset;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3127 0 0
2
5.90009e-315 5.39824e-315
0
12 Hex Display~
7 1081 239 0 16 19
10 25 24 23 96 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
559 0 0
2
5.90009e-315 5.40342e-315
0
9 Terminal~
194 1078 303 0 1 3
0 23
0
0 0 49520 180
4 ini3
7 -7 35 1
3 T87
-10 -32 11 -24
0
5 ini3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8488 0 0
2
5.90009e-315 5.4086e-315
0
9 Terminal~
194 1084 290 0 1 3
0 24
0
0 0 49520 180
4 ini2
7 -7 35 1
3 T88
-10 -32 11 -24
0
5 ini2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3392 0 0
2
5.90009e-315 5.41378e-315
0
9 Terminal~
194 1090 278 0 1 3
0 25
0
0 0 49520 180
4 ini1
7 -7 35 1
4 T124
-13 -32 15 -24
0
5 ini1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3952 0 0
2
5.90009e-315 5.41896e-315
0
9 Terminal~
194 1174 276 0 1 3
0 12
0
0 0 49520 180
4 qua1
7 -7 35 1
4 T126
-13 -32 15 -24
0
5 qua1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8186 0 0
2
5.90009e-315 5.42414e-315
0
9 Terminal~
194 1168 288 0 1 3
0 13
0
0 0 49520 180
4 qua2
7 -7 35 1
4 T127
-13 -32 15 -24
0
5 qua2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6571 0 0
2
5.90009e-315 5.42933e-315
0
9 Terminal~
194 1162 301 0 1 3
0 14
0
0 0 49520 180
4 qua3
7 -7 35 1
4 T128
-13 -32 15 -24
0
5 qua3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6167 0 0
2
5.90009e-315 5.43192e-315
0
12 Hex Display~
7 1165 237 0 16 19
10 12 13 14 2 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3566 0 0
2
5.90009e-315 5.43451e-315
0
9 Terminal~
194 912 133 0 1 3
0 26
0
0 0 49520 180
6 final2
-43 4 -1 12
4 T157
-13 -32 15 -24
0
7 final2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3371 0 0
2
5.90009e-315 5.4371e-315
0
12 Hex Display~
7 915 89 0 16 19
10 27 28 26 29 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP4
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4395 0 0
2
5.90009e-315 5.43969e-315
0
9 Terminal~
194 924 133 0 1 3
0 27
0
0 0 49520 180
6 final0
10 -11 52 -3
4 T156
-13 -32 15 -24
0
7 final0;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6822 0 0
2
5.90009e-315 5.44228e-315
0
9 Terminal~
194 918 133 0 1 3
0 28
0
0 0 49520 180
6 final1
6 5 48 13
4 T155
-13 -32 15 -24
0
7 final1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8953 0 0
2
5.90009e-315 5.44487e-315
0
9 Terminal~
194 906 133 0 1 3
0 29
0
0 0 49520 180
6 final3
-53 -9 -11 -1
4 T154
-13 -32 15 -24
0
7 final3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4635 0 0
2
5.90009e-315 5.44746e-315
0
9 Terminal~
194 985 774 0 1 3
0 18
0
0 0 49520 270
3 set
-17 6 4 14
3 T50
-10 -32 11 -24
0
4 set;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6596 0 0
2
5.90009e-315 5.45005e-315
0
2 +V
167 758 724 0 1 3
0 71
0
0 0 54256 0
2 5V
-7 -22 7 -14
3 V12
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3813 0 0
2
5.90009e-315 5.45264e-315
0
9 Inverter~
13 903 773 0 2 22
0 30 18
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
5639 0 0
2
5.90009e-315 5.45523e-315
0
9 Terminal~
194 918 733 0 1 3
0 30
0
0 0 49520 270
5 block
-31 -19 4 -11
3 T61
-10 -32 11 -24
0
6 block;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
429 0 0
2
5.90009e-315 5.45782e-315
0
7 Ground~
168 852 798 0 1 3
0 6
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5832 0 0
2
5.90009e-315 5.46041e-315
0
9 Terminal~
194 741 793 0 1 3
0 31
0
0 0 49520 90
6 clock3
-50 -5 -8 3
3 T22
-10 -32 11 -24
0
7 clock3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8856 0 0
2
5.90009e-315 5.463e-315
0
9 Terminal~
194 741 802 0 1 3
0 32
0
0 0 49520 90
6 clock2
-49 -5 -7 3
3 T21
-10 -32 11 -24
0
7 clock2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
469 0 0
2
5.90009e-315 5.46559e-315
0
9 Terminal~
194 741 766 0 1 3
0 33
0
0 0 49520 90
7 coluna3
-55 -7 -6 1
3 T20
-10 -32 11 -24
0
8 coluna3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4529 0 0
2
5.90009e-315 5.46818e-315
0
9 Terminal~
194 741 775 0 1 3
0 34
0
0 0 49520 90
7 coluna2
-55 -7 -6 1
3 T19
-10 -32 11 -24
0
8 coluna2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
88 0 0
2
5.90009e-315 5.47077e-315
0
9 Terminal~
194 741 784 0 1 3
0 35
0
0 0 49520 90
7 coluna1
-55 -7 -6 1
3 T18
-10 -32 11 -24
0
8 coluna1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3894 0 0
2
5.90009e-315 5.47207e-315
0
7 74LS153
119 806 791 0 14 29
0 71 33 34 35 31 32 97 98 99
100 6 101 30 102
0
0 0 4848 0
7 74LS153
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 512 1 0 0 0
1 U
6890 0 0
2
5.90009e-315 5.47336e-315
0
9 Terminal~
194 2624 620 0 1 3
0 27
0
0 0 49520 270
6 final0
-21 -15 21 -7
4 T161
-14 -32 14 -24
0
7 final0;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3257 0 0
2
5.90009e-315 5.47466e-315
0
9 Terminal~
194 2620 480 0 1 3
0 28
0
0 0 49520 270
6 final1
-21 -15 21 -7
4 T160
-14 -32 14 -24
0
7 final1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6612 0 0
2
5.90009e-315 5.47595e-315
0
9 Terminal~
194 2623 333 0 1 3
0 26
0
0 0 49520 270
6 final2
-21 -15 21 -7
4 T159
-14 -32 14 -24
0
7 final2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3556 0 0
2
5.90009e-315 5.47725e-315
0
9 Terminal~
194 2625 190 0 1 3
0 29
0
0 0 49520 270
6 final3
-21 -15 21 -7
4 T158
-14 -32 14 -24
0
7 final3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9143 0 0
2
5.90009e-315 5.47854e-315
0
9 Terminal~
194 1543 161 0 1 3
0 5
0
0 0 49520 90
7 letecla
-25 -15 24 -7
4 T150
-13 -32 15 -24
0
8 letecla;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8186 0 0
2
5.90009e-315 5.47984e-315
0
9 Inverter~
13 1583 159 0 2 22
0 5 73
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 11 0
1 U
3754 0 0
2
5.90009e-315 5.48113e-315
0
9 Terminal~
194 1676 70 0 1 3
0 18
0
0 0 49520 270
7 writeup
3 -5 52 3
4 T102
-13 -32 15 -24
0
8 writeup;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8708 0 0
2
5.90009e-315 5.48243e-315
0
9 Terminal~
194 1681 186 0 1 3
0 19
0
0 0 49520 270
6 readup
6 -5 48 3
4 T101
-13 -32 15 -24
0
7 readup;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3338 0 0
2
5.90009e-315 5.48372e-315
0
9 Terminal~
194 1681 154 0 1 3
0 19
0
0 0 49520 270
6 modoup
6 -5 48 3
3 T89
-10 -32 11 -24
0
7 modoup;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5546 0 0
2
5.90009e-315 5.48502e-315
0
9 2-In AND~
219 1638 168 0 3 22
0 73 36 19
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U23C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 13 0
1 U
3295 0 0
2
5.90009e-315 5.48631e-315
0
9 Terminal~
194 1598 215 0 1 3
0 36
0
0 0 49520 180
6 nvazio
3 -7 45 1
4 T147
-14 -32 14 -24
0
7 nvazio;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4923 0 0
2
5.90009e-315 5.48761e-315
0
9 Terminal~
194 2131 466 0 1 3
0 37
0
0 0 49520 270
7 output1
-25 -15 24 -7
3 T56
-11 -32 10 -24
0
8 output1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3248 0 0
2
5.90009e-315 5.4889e-315
0
9 Terminal~
194 2131 452 0 1 3
0 38
0
0 0 49520 270
7 output2
-25 -15 24 -7
3 T55
-11 -32 10 -24
0
8 output2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3139 0 0
2
5.90009e-315 5.4902e-315
0
9 Terminal~
194 2131 436 0 1 3
0 39
0
0 0 49520 270
7 output3
-25 -15 24 -7
3 T54
-11 -32 10 -24
0
8 output3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3285 0 0
2
5.90009e-315 5.49149e-315
0
9 Terminal~
194 2131 418 0 1 3
0 40
0
0 0 49520 270
7 output4
-25 -15 24 -7
3 T52
-11 -32 10 -24
0
8 output4;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
336 0 0
2
5.90009e-315 5.49279e-315
0
9 Terminal~
194 843 597 0 1 3
0 38
0
0 0 49520 270
7 output2
3 -7 52 1
3 T53
-10 -32 11 -24
0
8 output2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6582 0 0
2
5.90009e-315 5.49408e-315
0
9 Terminal~
194 843 615 0 1 3
0 37
0
0 0 49520 270
7 output1
3 -7 52 1
3 T51
-10 -32 11 -24
0
8 output1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3546 0 0
2
5.90009e-315 5.49538e-315
0
9 Terminal~
194 843 579 0 1 3
0 39
0
0 0 49520 270
7 output3
3 -7 52 1
3 T49
-10 -32 11 -24
0
8 output3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
893 0 0
2
5.90009e-315 5.49667e-315
0
9 Terminal~
194 843 561 0 1 3
0 40
0
0 0 49520 270
7 output4
3 -7 52 1
3 T48
-10 -32 11 -24
0
8 output4;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8998 0 0
2
5.90009e-315 5.49797e-315
0
9 Terminal~
194 1791 1554 0 1 3
0 36
0
0 0 49520 270
6 nvazio
-13 -14 29 -6
4 T149
-14 -32 14 -24
0
7 nvazio;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5979 0 0
2
5.90009e-315 5.49926e-315
0
9 Terminal~
194 2274 188 0 1 3
0 20
0
0 0 49520 90
4 modo
-40 -7 -12 1
4 T145
-14 -32 14 -24
0
5 modo;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3835 0 0
2
44521.8 33
0
9 Terminal~
194 2273 179 0 1 3
0 41
0
0 0 49520 90
5 psave
-41 -12 -6 -4
4 T139
-14 -32 14 -24
0
6 psave;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
750 0 0
2
44521.8 34
0
5 7415~
219 2361 186 0 4 22
0 41 20 7 21
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U26A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 16 0
1 U
849 0 0
2
44521.8 35
0
9 Terminal~
194 2474 621 0 1 3
0 42
0
0 0 49520 90
4 reg0
-14 -15 14 -7
4 T143
-14 -32 14 -24
0
5 reg0;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4693 0 0
2
44521.8 36
0
9 Terminal~
194 2477 481 0 1 3
0 43
0
0 0 49520 90
4 reg1
-14 -15 14 -7
4 T142
-14 -32 14 -24
0
5 reg1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4775 0 0
2
44521.8 37
0
9 Terminal~
194 2473 333 0 1 3
0 44
0
0 0 49520 90
4 reg2
-14 -15 14 -7
4 T141
-14 -32 14 -24
0
5 reg2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9572 0 0
2
44521.8 38
0
9 Terminal~
194 2476 191 0 1 3
0 45
0
0 0 49520 90
4 reg3
-14 -15 14 -7
4 T140
-14 -32 14 -24
0
5 reg3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3761 0 0
2
44521.8 39
0
9 Terminal~
194 1891 482 0 1 3
0 41
0
0 0 49520 270
5 psave
-18 -15 17 -7
4 T138
-14 -32 14 -24
0
6 psave;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6765 0 0
2
44521.8 40
0
9 Terminal~
194 1892 536 0 1 3
0 43
0
0 0 49520 270
4 reg1
-15 -15 13 -7
4 T137
-14 -32 14 -24
0
5 reg1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7938 0 0
2
44521.8 41
0
9 Terminal~
194 1892 551 0 1 3
0 42
0
0 0 49520 270
4 reg0
-15 -15 13 -7
4 T136
-14 -32 14 -24
0
5 reg0;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
55 0 0
2
44521.8 42
0
9 Terminal~
194 1892 520 0 1 3
0 44
0
0 0 49520 270
4 reg2
-15 -15 13 -7
4 T117
-14 -32 14 -24
0
5 reg2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5610 0 0
2
44521.8 43
0
9 Terminal~
194 1892 505 0 1 3
0 45
0
0 0 49520 270
4 reg3
-15 -15 13 -7
4 T116
-14 -32 14 -24
0
5 reg3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3322 0 0
2
44521.8 44
0
9 Terminal~
194 2049 1254 0 1 3
0 20
0
0 0 49520 0
4 modo
-14 -22 14 -14
3 T76
-11 -32 10 -24
0
5 modo;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5914 0 0
2
44521.8 45
0
9 Terminal~
194 1901 1272 0 1 3
0 19
0
0 0 49520 0
6 modoup
-50 -6 -8 2
3 T72
-11 -32 10 -24
0
7 modoup;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8748 0 0
2
44521.8 46
0
5 4013~
219 1967 1300 0 6 22
0 6 74 19 8 103 20
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U15A
21 -54 49 -46
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 15 0
1 U
5830 0 0
2
44521.8 47
0
9 Terminal~
194 1967 1333 0 1 3
0 8
0
0 0 49520 180
6 mododw
7 -7 49 1
3 T66
-11 -32 10 -24
0
7 mododw;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9153 0 0
2
44521.8 48
0
2 +V
167 1920 1240 0 1 3
0 74
0
0 0 54256 0
2 5V
-7 -22 7 -14
3 V14
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9220 0 0
2
44521.8 49
0
7 Ground~
168 1936 1326 0 1 3
0 6
0
0 0 53360 0
0
5 GND22
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7901 0 0
2
44521.8 50
0
2 +V
167 2026 268 0 1 3
0 75
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4571 0 0
2
44521.8 51
0
7 Ground~
168 1679 1321 0 1 3
0 6
0
0 0 53360 0
0
5 GND20
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7796 0 0
2
5.90009e-315 5.50056e-315
0
2 +V
167 1663 1235 0 1 3
0 76
0
0 0 54256 0
2 5V
-7 -22 7 -14
3 V11
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3907 0 0
2
5.90009e-315 5.50185e-315
0
9 Terminal~
194 1710 1328 0 1 3
0 46
0
0 0 49520 180
6 dddown
7 -7 49 1
3 T65
-11 -32 10 -24
0
7 dddown;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4389 0 0
2
5.90009e-315 5.50315e-315
0
2 +V
167 1293 946 0 1 3
0 77
0
0 0 54256 0
2 5V
-7 -22 7 -14
3 V10
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7762 0 0
2
5.90009e-315 5.50444e-315
0
7 74LS191
135 1641 1024 0 14 29
0 6 15 22 20 6 6 6 6 104
105 2 14 13 12
0
0 0 4848 0
7 74LS191
-24 -51 25 -43
3 U25
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
6723 0 0
2
5.90009e-315 5.50574e-315
0
9 Terminal~
194 1699 1043 0 1 3
0 14
0
0 0 49520 270
4 qua3
6 -7 34 1
4 T130
-13 -32 15 -24
0
5 qua3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6871 0 0
2
5.90009e-315 5.50703e-315
0
9 Terminal~
194 1699 1052 0 1 3
0 13
0
0 0 49520 270
4 qua2
6 -7 34 1
4 T131
-13 -32 15 -24
0
5 qua2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4198 0 0
2
5.90009e-315 5.50833e-315
0
9 Terminal~
194 1699 1061 0 1 3
0 12
0
0 0 49520 270
4 qua1
5 -6 33 2
4 T132
-13 -32 15 -24
0
5 qua1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
970 0 0
2
5.90009e-315 5.50963e-315
0
9 Terminal~
194 1739 1024 0 1 3
0 2
0
0 0 49520 0
5 qoito
-17 -22 18 -14
4 T133
-14 -32 14 -24
0
6 qoito;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
319 0 0
2
5.90009e-315 5.51092e-315
0
7 Ground~
168 1592 1117 0 1 3
0 6
0
0 0 53360 0
0
5 GND24
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3663 0 0
2
5.90009e-315 5.51222e-315
0
9 Terminal~
194 1567 1026 0 1 3
0 20
0
0 0 49520 90
4 modo
-35 -6 -7 2
4 T134
-14 -32 14 -24
0
5 modo;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3512 0 0
2
5.90009e-315 5.51286e-315
0
9 Terminal~
194 1567 1008 0 1 3
0 15
0
0 0 49520 90
2 pq
-28 -5 -14 3
4 T135
-14 -32 14 -24
0
3 pq;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7555 0 0
2
5.90009e-315 5.51351e-315
0
9 Terminal~
194 1774 155 0 1 3
0 20
0
0 0 49520 270
4 modo
6 -5 34 3
4 T104
-13 -32 15 -24
0
5 modo;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9776 0 0
2
5.90009e-315 5.51416e-315
0
9 Terminal~
194 1678 1460 0 1 3
0 20
0
0 0 49520 90
4 modo
-38 -6 -10 2
3 T84
-11 -32 10 -24
0
5 modo;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6596 0 0
2
5.90009e-315 5.51481e-315
0
9 2-In AND~
219 1736 1467 0 3 22
0 20 7 46
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U23A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
6750 0 0
2
5.90009e-315 5.51545e-315
0
9 Terminal~
194 1679 1478 0 1 3
0 7
0
0 0 49520 90
5 wrout
-41 -6 -6 2
4 T122
-14 -32 14 -24
0
6 wrout;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9636 0 0
2
5.90009e-315 5.5161e-315
0
9 Terminal~
194 1807 1468 0 1 3
0 46
0
0 0 49520 270
6 dddown
-21 -15 21 -7
4 T123
-14 -32 14 -24
0
7 dddown;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5369 0 0
2
5.90009e-315 5.51675e-315
0
9 Terminal~
194 1808 1524 0 1 3
0 47
0
0 0 49520 270
4 ddup
-15 -15 13 -7
4 T121
-14 -32 14 -24
0
5 ddup;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8555 0 0
2
5.90009e-315 5.5174e-315
0
9 2-In AND~
219 1737 1523 0 3 22
0 48 36 47
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U23B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 13 0
1 U
4690 0 0
2
5.90009e-315 5.51804e-315
0
9 Terminal~
194 1679 1516 0 1 3
0 48
0
0 0 49520 90
6 nclock
-45 -6 -3 2
4 T125
-14 -32 14 -24
0
7 nclock;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9145 0 0
2
5.90009e-315 5.51869e-315
0
9 Terminal~
194 1294 746 0 1 3
0 2
0
0 0 49520 180
5 qoito
-13 11 22 19
3 T90
-10 -32 11 -24
0
6 qoito;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5246 0 0
2
5.90009e-315 5.51934e-315
0
9 Terminal~
194 1276 745 0 1 3
0 14
0
0 0 49520 180
4 qua3
-20 1 8 9
3 T86
-10 -32 11 -24
0
5 qua3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9111 0 0
2
5.90009e-315 5.51999e-315
0
8 2-In OR~
219 1282 695 0 3 22
0 14 2 80
0
0 0 624 90
6 74LS32
-21 -24 21 -16
4 U19C
29 -3 57 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
6717 0 0
2
5.90009e-315 5.52063e-315
0
9 2-In AND~
219 1277 628 0 3 22
0 79 80 78
0
0 0 624 90
6 74LS08
-21 -24 21 -16
4 U20D
17 -5 45 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 10 0
1 U
3487 0 0
2
5.90009e-315 5.52128e-315
0
9 Inverter~
13 1411 962 0 2 22
0 82 81
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U3B
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 11 0
1 U
9604 0 0
2
5.90009e-315 5.52193e-315
0
9 Terminal~
194 1232 1674 0 1 3
0 8
0
0 0 49520 270
7 pinicio
-25 -15 24 -7
3 T85
-11 -32 10 -24
0
8 pinicio;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3921 0 0
2
5.90009e-315 5.52258e-315
0
9 Terminal~
194 1036 1684 0 1 3
0 20
0
0 0 49520 90
4 modo
-36 -6 -8 2
4 T105
-14 -32 14 -24
0
5 modo;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8146 0 0
2
5.90009e-315 5.52322e-315
0
5 4081~
219 1147 1673 0 3 22
0 16 20 8
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U22B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 12 0
1 U
4506 0 0
2
5.90009e-315 5.52387e-315
0
9 Terminal~
194 1034 1618 0 1 3
0 7
0
0 0 49520 90
5 wrout
-39 -6 -4 2
4 T112
-14 -32 14 -24
0
6 wrout;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5386 0 0
2
5.90009e-315 5.52452e-315
0
5 4081~
219 1085 1625 0 3 22
0 7 48 16
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U22A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 12 0
1 U
7847 0 0
2
5.90009e-315 5.52517e-315
0
9 Terminal~
194 1034 1636 0 1 3
0 48
0
0 0 49520 90
6 nclock
-43 -5 -1 3
4 T113
-14 -32 14 -24
0
7 nclock;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9261 0 0
2
5.90009e-315 5.52581e-315
0
9 Terminal~
194 233 664 0 1 3
0 49
0
0 0 49520 270
7 clinha4
3 -4 52 4
4 T111
-14 -32 14 -24
0
8 clinha4;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8231 0 0
2
5.90009e-315 5.52646e-315
0
9 Terminal~
194 233 673 0 1 3
0 50
0
0 0 49520 270
7 clinha3
1 -4 50 4
4 T110
-14 -32 14 -24
0
8 clinha3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3756 0 0
2
5.90009e-315 5.52711e-315
0
9 Terminal~
194 233 691 0 1 3
0 51
0
0 0 49520 270
7 clinha1
2 -4 51 4
4 T109
-14 -32 14 -24
0
8 clinha1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6760 0 0
2
5.90009e-315 5.52776e-315
0
9 Terminal~
194 233 682 0 1 3
0 52
0
0 0 49520 270
7 clinha2
2 -4 51 4
4 T108
-14 -32 14 -24
0
8 clinha2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
351 0 0
2
5.90009e-315 5.52841e-315
0
9 Terminal~
194 96 674 0 1 3
0 53
0
0 0 49520 90
6 clock1
-45 -6 -3 2
4 T107
-14 -32 14 -24
0
7 clock1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5352 0 0
2
5.90009e-315 5.52905e-315
0
9 Terminal~
194 96 683 0 1 3
0 54
0
0 0 49520 90
6 clock0
-48 -4 -6 4
4 T106
-14 -32 14 -24
0
7 clock0;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
485 0 0
2
5.90009e-315 5.5297e-315
0
7 74LS139
118 181 654 0 14 29
0 53 54 6 53 54 6 62 65 64
63 49 50 52 51
0
0 0 13040 0
7 74LS139
-24 -51 25 -43
3 U21
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
113 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+[%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
13 type: digital
5 DIP16
29

0 3 2 1 13 14 15 7 6 5
4 9 10 11 12 3 2 1 13 14
15 7 6 5 4 9 10 11 12 70
65 0 0 0 1 1 0 0
1 U
452 0 0
2
5.90009e-315 5.53035e-315
0
7 74LS293
154 191 540 0 8 17
0 6 6 92 54 31 32 53 54
0
0 0 4848 0
7 74LS293
-24 -35 25 -27
2 U1
-7 -36 7 -28
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 0 1 0 0 0
1 U
643 0 0
2
5.90009e-315 5.531e-315
0
9 Terminal~
194 1164 658 0 1 3
0 20
0
0 0 49520 90
4 modo
-32 -6 -4 2
3 T92
-10 -32 11 -24
0
5 modo;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5563 0 0
2
44521.8 52
0
8 2-In OR~
219 1346 694 0 3 22
0 13 2 84
0
0 0 624 90
6 74LS32
-21 -24 21 -16
4 U19A
29 -3 57 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
934 0 0
2
44521.8 53
0
9 2-In AND~
219 1341 628 0 3 22
0 79 84 85
0
0 0 624 90
6 74LS08
-21 -24 21 -16
4 U20A
17 -5 45 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
3240 0 0
2
44521.8 54
0
9 Inverter~
13 1221 656 0 2 22
0 20 79
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
3233 0 0
2
44521.8 55
0
9 Terminal~
194 1340 741 0 1 3
0 13
0
0 0 49520 180
4 qua2
-20 1 8 9
3 T91
-10 -32 11 -24
0
5 qua2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3635 0 0
2
44521.8 56
0
9 Terminal~
194 1358 741 0 1 3
0 2
0
0 0 49520 180
5 qoito
-12 11 23 19
3 T93
-10 -32 11 -24
0
6 qoito;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3547 0 0
2
44521.8 57
0
9 2-In AND~
219 1413 630 0 3 22
0 79 83 86
0
0 0 624 90
6 74LS08
-21 -24 21 -16
4 U20B
17 -5 45 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
483 0 0
2
44521.8 58
0
8 2-In OR~
219 1418 696 0 3 22
0 12 2 83
0
0 0 624 90
6 74LS32
-21 -24 21 -16
4 U19B
29 -3 57 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
6126 0 0
2
44521.8 59
0
9 Terminal~
194 1412 743 0 1 3
0 12
0
0 0 49520 180
4 qua1
-20 1 8 9
3 T95
-10 -32 11 -24
0
5 qua1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7368 0 0
2
44521.8 60
0
9 Terminal~
194 1430 743 0 1 3
0 2
0
0 0 49520 180
5 qoito
-13 11 22 19
4 T103
-13 -32 15 -24
0
6 qoito;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3925 0 0
2
44521.8 61
0
9 Terminal~
194 1431 1044 0 1 3
0 23
0
0 0 49520 270
4 ini3
6 -6 34 2
3 T98
-10 -32 11 -24
0
5 ini3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6187 0 0
2
44521.8 62
0
9 Terminal~
194 1431 1053 0 1 3
0 24
0
0 0 49520 270
4 ini2
6 -7 34 1
3 T99
-10 -32 11 -24
0
5 ini2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5866 0 0
2
44521.8 63
0
9 Terminal~
194 1431 1062 0 1 3
0 25
0
0 0 49520 270
4 ini1
5 -6 33 2
4 T100
-13 -32 15 -24
0
5 ini1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6650 0 0
2
44521.8 64
0
9 Terminal~
194 1447 523 0 1 3
0 23
0
0 0 49520 90
4 ini3
-32 -6 -4 2
3 T97
-10 -32 11 -24
0
5 ini3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8814 0 0
2
44521.8 65
0
9 Terminal~
194 1447 532 0 1 3
0 24
0
0 0 49520 90
4 ini2
-32 -6 -4 2
3 T96
-10 -32 11 -24
0
5 ini2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4714 0 0
2
44521.8 66
0
9 Terminal~
194 1447 541 0 1 3
0 25
0
0 0 49520 90
4 ini1
-32 -6 -4 2
3 T94
-10 -32 11 -24
0
5 ini1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9875 0 0
2
44521.8 67
0
6 74LS83
105 1523 548 0 14 29
0 6 23 24 25 6 78 85 86 6
106 9 10 11 6
0
0 0 4848 0
6 74LS83
-21 -60 21 -52
3 U16
-10 -61 11 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
8220 0 0
2
44521.8 68
0
7 Ground~
168 1475 664 0 1 3
0 6
0
0 0 53360 0
0
5 GND25
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3691 0 0
2
44521.8 69
0
9 2-In AND~
219 1082 1495 0 3 22
0 17 2 56
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
5196 0 0
2
44521.8 70
0
9 2-In AND~
219 1387 1495 0 3 22
0 48 87 55
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
6182 0 0
2
44521.8 71
0
9 Terminal~
194 166 486 0 1 3
0 48
0
0 0 49520 270
6 nclock
2 -4 44 4
3 T83
-10 -32 11 -24
0
7 nclock;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6326 0 0
2
44521.8 72
0
9 Inverter~
13 1326 1504 0 2 22
0 2 87
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
3247 0 0
2
44521.8 73
0
9 Terminal~
194 1452 1486 0 1 3
0 55
0
0 0 49520 0
6 ordown
-21 -22 21 -14
3 T82
-11 -32 10 -24
0
7 ordown;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5235 0 0
2
44521.8 74
0
9 Terminal~
194 1267 1493 0 1 3
0 2
0
0 0 49520 0
5 qoito
-17 -22 18 -14
3 T81
-11 -32 10 -24
0
6 qoito;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9260 0 0
2
44521.8 75
0
9 Terminal~
194 1304 1477 0 1 3
0 48
0
0 0 49520 0
6 nclock
-20 -22 22 -14
3 T80
-11 -32 10 -24
0
7 nclock;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
583 0 0
2
44521.8 76
0
9 Terminal~
194 1000 1477 0 1 3
0 17
0
0 0 49520 0
5 clock
-17 -22 18 -14
3 T77
-11 -32 10 -24
0
6 clock;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3471 0 0
2
44521.8 77
0
9 Terminal~
194 1035 1494 0 1 3
0 2
0
0 0 49520 0
5 qoito
-17 -22 18 -14
3 T78
-11 -32 10 -24
0
6 qoito;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7124 0 0
2
44521.8 78
0
9 Terminal~
194 1134 1486 0 1 3
0 56
0
0 0 49520 0
4 orup
-14 -22 14 -14
3 T79
-11 -32 10 -24
0
5 orup;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6160 0 0
2
44521.8 79
0
5 4013~
219 1710 1295 0 6 22
0 6 76 47 46 107 3
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U18B
21 -54 49 -46
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 9 0
1 U
4732 0 0
2
44521.8 80
0
9 Terminal~
194 1644 1267 0 1 3
0 47
0
0 0 49520 0
4 ddup
-14 -21 14 -13
3 T71
-11 -32 10 -24
0
5 ddup;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8836 0 0
2
44521.8 81
0
9 Terminal~
194 1792 1249 0 1 3
0 3
0
0 0 49520 0
5 ddout
-17 -22 18 -14
3 T70
-11 -32 10 -24
0
6 ddout;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3346 0 0
2
44521.8 82
0
5 4013~
219 1400 1295 0 6 22
0 6 88 56 55 108 4
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U18A
21 -54 49 -46
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 9 0
1 U
8546 0 0
2
44521.8 83
0
2 +V
167 1339 1247 0 1 3
0 88
0
0 0 54256 0
3 10V
-11 -22 10 -14
3 V17
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8607 0 0
2
44521.8 84
0
9 Terminal~
194 1299 1266 0 1 3
0 56
0
0 0 49520 0
4 orup
-14 -22 14 -14
3 T69
-11 -32 10 -24
0
5 orup;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5781 0 0
2
44521.8 85
0
9 Terminal~
194 1332 1304 0 1 3
0 55
0
0 0 49520 0
6 ordown
-21 -22 21 -14
3 T68
-11 -32 10 -24
0
7 ordown;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6991 0 0
2
44521.8 86
0
9 Terminal~
194 1482 1249 0 1 3
0 4
0
0 0 49520 0
5 orout
-17 -22 18 -14
3 T67
-11 -32 10 -24
0
6 orout;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9631 0 0
2
44521.8 87
0
7 Ground~
168 1371 1337 0 1 3
0 6
0
0 0 53360 0
0
5 GND21
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8381 0 0
2
44521.8 88
0
7 Ground~
168 1076 1338 0 1 3
0 6
0
0 0 53360 0
0
5 GND23
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6697 0 0
2
44521.8 89
0
9 Terminal~
194 1187 1250 0 1 3
0 7
0
0 0 49520 0
5 wrout
-17 -22 18 -14
3 T75
-11 -32 10 -24
0
6 wrout;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3463 0 0
2
44521.8 90
0
9 Terminal~
194 1037 1305 0 1 3
0 16
0
0 0 49520 0
6 wrdown
-21 -22 21 -14
3 T74
-11 -32 10 -24
0
7 wrdown;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9605 0 0
2
44521.8 91
0
2 +V
167 1044 1248 0 1 3
0 90
0
0 0 54256 0
3 10V
-11 -22 10 -14
3 V16
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
936 0 0
2
44521.8 92
0
5 4013~
219 1105 1296 0 6 22
0 6 90 89 16 109 7
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U17B
21 -54 49 -46
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 8 0
1 U
9813 0 0
2
44521.8 93
0
7 74LS193
137 1374 1025 0 14 29
0 8 77 81 6 6 6 6 6 110
111 82 23 24 25
0
0 0 4848 0
7 74LS193
-24 -51 25 -43
3 U14
-11 -52 10 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
5286 0 0
2
44521.8 94
0
7 Ground~
168 1325 1113 0 1 3
0 6
0
0 0 53360 0
0
5 GND19
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9179 0 0
2
44521.8 95
0
9 Terminal~
194 1260 989 0 1 3
0 8
0
0 0 49520 0
7 pinicio
-25 -22 24 -14
3 T63
-11 -32 10 -24
0
8 pinicio;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3718 0 0
2
44521.8 96
0
7 Ground~
168 1904 302 0 1 3
0 6
0
0 0 53360 0
0
5 GND18
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4375 0 0
2
5.90009e-315 5.53164e-315
0
5 4013~
219 2541 225 0 6 22
0 6 45 21 6 112 29
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U10A
23 -61 51 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 5 0
1 U
3616 0 0
2
5.90009e-315 5.53229e-315
0
7 Ground~
168 2647 149 0 1 3
0 6
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7808 0 0
2
5.90009e-315 5.53294e-315
0
7 Ground~
168 2541 249 0 1 3
0 6
0
0 0 53360 0
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7498 0 0
2
5.90009e-315 5.53359e-315
0
7 Ground~
168 2538 393 0 1 3
0 6
0
0 0 53360 0
0
5 GND11
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9736 0 0
2
5.90009e-315 5.53423e-315
0
7 Ground~
168 2645 290 0 1 3
0 6
0
0 0 53360 0
0
5 GND12
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9454 0 0
2
5.90009e-315 5.53488e-315
0
5 4013~
219 2538 367 0 6 22
0 6 44 21 6 113 26
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U10B
23 -61 51 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 5 0
1 U
4639 0 0
2
5.90009e-315 5.53553e-315
0
7 Ground~
168 2538 539 0 1 3
0 6
0
0 0 53360 0
0
5 GND13
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3831 0 0
2
5.90009e-315 5.53618e-315
0
7 Ground~
168 2645 434 0 1 3
0 6
0
0 0 53360 0
0
5 GND14
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3538 0 0
2
5.90009e-315 5.53682e-315
0
5 4013~
219 2538 515 0 6 22
0 6 43 21 6 114 28
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U11A
23 -61 51 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 6 0
1 U
5949 0 0
2
5.90009e-315 5.53747e-315
0
7 Ground~
168 2541 679 0 1 3
0 6
0
0 0 53360 0
0
5 GND15
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7130 0 0
2
5.90009e-315 5.53812e-315
0
7 Ground~
168 2641 578 0 1 3
0 6
0
0 0 53360 0
0
5 GND16
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4115 0 0
2
5.90009e-315 5.53877e-315
0
5 4013~
219 2541 655 0 6 22
0 6 42 21 6 115 27
0
0 0 4720 0
4 4013
10 -60 38 -52
4 U11B
23 -61 51 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 6 0
1 U
3197 0 0
2
5.90009e-315 5.53941e-315
0
7 74LS245
64 1959 312 0 18 37
0 116 117 118 41 45 44 43 42 119
120 121 75 40 39 38 37 6 20
0
0 0 4848 0
7 74LS245
-24 -60 25 -52
3 U13
-11 -61 10 -53
0
16 DVCC=20;DGND=10;
192 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i]
+ [%20bi %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP14
37

0 9 8 7 6 5 4 3 2 11
12 13 14 15 16 17 18 19 1 9
8 7 6 5 4 3 2 11 12 13
14 15 16 17 18 19 1 0
65 0 0 512 1 0 0 0
1 U
813 0 0
2
5.90009e-315 5.54006e-315
0
7 Ground~
168 1624 479 0 1 3
0 6
0
0 0 53360 0
0
5 GND17
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3396 0 0
2
5.90009e-315 5.54071e-315
0
6 1K RAM
79 1672 404 0 20 41
0 6 6 6 6 6 6 6 9 10
11 122 123 124 41 45 44 43 42 66
20
0
0 0 4848 0
5 RAM1K
-17 -19 18 -11
3 U12
-11 -70 10 -62
0
16 DVCC=22;DGND=11;
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 512 1 0 0 0
1 U
6348 0 0
2
5.90009e-315 5.54136e-315
0
6 74LS83
105 547 569 0 14 29
0 6 6 31 32 6 51 91 52 6
57 58 60 59 125
0
0 0 4848 0
6 74LS83
-21 -60 21 -52
2 U4
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
583 0 0
2
44521.8 97
0
9 Inverter~
13 420 587 0 2 22
0 50 91
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
922 0 0
2
44521.8 98
0
9 Terminal~
194 489 580 0 1 3
0 51
0
0 0 49520 90
7 clinha1
-55 -7 -6 1
3 T23
-10 -32 11 -24
0
8 clinha1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4442 0 0
2
44521.8 99
0
9 Terminal~
194 393 589 0 1 3
0 50
0
0 0 49520 90
7 clinha3
-55 -7 -6 1
3 T24
-10 -32 11 -24
0
8 clinha3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5893 0 0
2
44521.8 100
0
9 Terminal~
194 489 598 0 1 3
0 52
0
0 0 49520 90
7 clinha2
-55 -7 -6 1
3 T25
-10 -32 11 -24
0
8 clinha2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3814 0 0
2
44521.8 101
0
7 Ground~
168 506 635 0 1 3
0 6
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3637 0 0
2
44521.8 102
0
9 Terminal~
194 483 562 0 1 3
0 32
0
0 0 49520 90
6 clock2
-48 -6 -6 2
3 T26
-10 -32 11 -24
0
7 clock2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6890 0 0
2
44521.8 103
0
9 Terminal~
194 616 561 0 1 3
0 57
0
0 0 49520 270
3 sn3
12 -4 33 4
3 T30
-10 -32 11 -24
0
4 sn3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3933 0 0
2
44521.8 104
0
9 Terminal~
194 616 570 0 1 3
0 58
0
0 0 49520 270
3 sn2
12 -4 33 4
3 T31
-10 -32 11 -24
0
4 sn2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3432 0 0
2
44521.8 105
0
9 Terminal~
194 616 588 0 1 3
0 59
0
0 0 49520 270
3 sn0
12 -4 33 4
3 T32
-10 -32 11 -24
0
4 sn0;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3704 0 0
2
44521.8 106
0
9 Terminal~
194 616 579 0 1 3
0 60
0
0 0 49520 270
3 sn1
12 -4 33 4
3 T33
-10 -32 11 -24
0
4 sn1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9222 0 0
2
44521.8 107
0
9 Terminal~
194 483 553 0 1 3
0 31
0
0 0 49520 90
6 clock3
-48 -6 -6 2
3 T27
-10 -32 11 -24
0
7 clock3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8831 0 0
2
44521.8 108
0
9 Terminal~
194 483 723 0 1 3
0 32
0
0 0 49520 90
6 clock2
-48 -6 -6 2
3 T38
-10 -32 11 -24
0
7 clock2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9689 0 0
2
44521.8 109
0
9 Inverter~
13 516 721 0 2 22
0 32 61
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
469 0 0
2
44521.8 110
0
9 Terminal~
194 584 713 0 1 3
0 61
0
0 0 49520 270
3 se3
12 -4 33 4
3 T37
-10 -32 11 -24
0
4 se3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3309 0 0
2
44521.8 111
0
9 Terminal~
194 584 722 0 1 3
0 61
0
0 0 49520 270
3 se2
12 -4 33 4
3 T36
-10 -32 11 -24
0
4 se2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4792 0 0
2
44521.8 112
0
9 Terminal~
194 584 740 0 1 3
0 31
0
0 0 49520 270
3 se0
12 -4 33 4
3 T35
-10 -32 11 -24
0
4 se0;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3834 0 0
2
44521.8 113
0
9 Terminal~
194 584 731 0 1 3
0 61
0
0 0 49520 270
3 se1
12 -4 33 4
3 T34
-10 -32 11 -24
0
4 se1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5683 0 0
2
44521.8 114
0
9 Terminal~
194 535 741 0 1 3
0 31
0
0 0 49520 90
6 clock3
-48 -6 -6 2
3 T29
-10 -32 11 -24
0
7 clock3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5248 0 0
2
44521.8 115
0
9 Terminal~
194 166 466 0 1 3
0 17
0
0 0 49520 270
5 clock
5 -4 40 4
3 T28
-10 -32 11 -24
0
6 clock;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7816 0 0
2
44521.8 116
0
9 2-In AND~
219 105 549 0 3 22
0 17 30 92
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3496 0 0
2
44521.8 117
0
9 Terminal~
194 58 560 0 1 3
0 30
0
0 0 49520 90
5 block
-18 -15 17 -7
3 T62
-10 -32 11 -24
0
6 block;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3615 0 0
2
44521.8 118
0
9 Terminal~
194 741 544 0 1 3
0 62
0
0 0 49520 90
6 linha4
-47 -15 -5 -7
3 T47
-10 -32 11 -24
0
7 linha4;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7894 0 0
2
44521.8 119
0
9 Terminal~
194 741 616 0 1 3
0 31
0
0 0 49520 90
3 se0
-34 -6 -13 2
3 T46
-10 -32 11 -24
0
4 se0;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7766 0 0
2
44521.8 120
0
9 Terminal~
194 741 607 0 1 3
0 59
0
0 0 49520 90
3 sn0
-34 -6 -13 2
3 T45
-10 -32 11 -24
0
4 sn0;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9666 0 0
2
44521.8 121
0
9 Terminal~
194 741 598 0 1 3
0 61
0
0 0 49520 90
3 se1
-35 -6 -14 2
3 T44
-10 -32 11 -24
0
4 se1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8160 0 0
2
44521.8 122
0
9 Terminal~
194 741 589 0 1 3
0 60
0
0 0 49520 90
3 sn1
-35 -6 -14 2
3 T43
-10 -32 11 -24
0
4 sn1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5699 0 0
2
44521.8 123
0
9 Terminal~
194 741 580 0 1 3
0 61
0
0 0 49520 90
3 se2
-36 -5 -15 3
3 T42
-10 -32 11 -24
0
4 se2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9122 0 0
2
44521.8 124
0
9 Terminal~
194 741 571 0 1 3
0 58
0
0 0 49520 90
3 sn2
-35 -6 -14 2
3 T41
-10 -32 11 -24
0
4 sn2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8786 0 0
2
44521.8 125
0
9 Terminal~
194 741 562 0 1 3
0 61
0
0 0 49520 90
3 se3
-36 -6 -15 2
3 T40
-10 -32 11 -24
0
4 se3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8644 0 0
2
44521.8 126
0
9 Terminal~
194 741 553 0 1 3
0 57
0
0 0 49520 90
3 sn3
-35 -6 -14 2
3 T39
-10 -32 11 -24
0
4 sn3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3439 0 0
2
44521.8 127
0
7 Ground~
168 739 645 0 1 3
0 6
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3241 0 0
2
44521.8 128
0
7 74LS157
122 784 578 0 14 29
0 62 57 61 58 61 60 61 59 31
6 40 39 38 37
0
0 0 4848 0
7 74LS157
-24 -60 25 -52
2 U6
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
8130 0 0
2
44521.8 129
0
9 Terminal~
194 514 366 0 1 3
0 33
0
0 0 49520 180
7 coluna3
4 -7 53 1
3 T17
-10 -32 11 -24
0
8 coluna3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5945 0 0
2
44521.8 130
0
9 Terminal~
194 433 368 0 1 3
0 34
0
0 0 49520 180
7 coluna2
4 -7 53 1
3 T16
-10 -32 11 -24
0
8 coluna2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4456 0 0
2
44521.8 131
0
9 Terminal~
194 343 403 0 1 3
0 35
0
0 0 49520 180
7 coluna1
4 -7 53 1
3 T15
-10 -32 11 -24
0
8 coluna1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5515 0 0
2
44521.8 132
0
9 Terminal~
194 282 532 0 1 3
0 31
0
0 0 49520 270
6 clock3
2 -4 44 4
3 T14
-10 -32 11 -24
0
7 clock3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3289 0 0
2
44521.8 133
0
9 Terminal~
194 282 541 0 1 3
0 32
0
0 0 49520 270
6 clock2
2 -5 44 3
3 T13
-10 -32 11 -24
0
7 clock2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8691 0 0
2
44521.8 134
0
2 +V
167 343 55 0 1 3
0 93
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9388 0 0
2
44521.8 135
0
9 Terminal~
194 206 155 0 1 3
0 63
0
0 0 49520 90
6 linha1
-12 -17 30 -9
3 T12
-10 -32 11 -24
0
7 linha1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7836 0 0
2
44521.8 136
0
9 Terminal~
194 206 218 0 1 3
0 64
0
0 0 49520 90
6 linha2
-21 -15 21 -7
3 T11
-10 -32 11 -24
0
7 linha2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8355 0 0
2
44521.8 137
0
9 Terminal~
194 204 281 0 1 3
0 65
0
0 0 49520 90
6 linha3
-21 -15 21 -7
3 T10
-10 -32 11 -24
0
7 linha3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3374 0 0
2
44521.8 138
0
9 Terminal~
194 205 344 0 1 3
0 62
0
0 0 49520 90
6 linha4
-21 -15 21 -7
2 T9
-7 -32 7 -24
0
7 linha4;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9602 0 0
2
44521.8 139
0
9 Terminal~
194 233 646 0 1 3
0 64
0
0 0 49520 270
6 linha2
2 -5 44 3
2 T8
-7 -32 7 -24
0
7 linha2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3548 0 0
2
44521.8 140
0
9 Terminal~
194 233 655 0 1 3
0 63
0
0 0 49520 270
6 linha1
2 -4 44 4
2 T7
-7 -32 7 -24
0
7 linha1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3407 0 0
2
44521.8 141
0
9 Terminal~
194 233 637 0 1 3
0 65
0
0 0 49520 270
6 linha3
2 -4 44 4
2 T6
-7 -32 7 -24
0
7 linha3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3554 0 0
2
44521.8 142
0
9 Terminal~
194 233 628 0 1 3
0 62
0
0 0 49520 270
6 linha4
2 -4 44 4
2 T5
-7 -32 7 -24
0
7 linha4;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8535 0 0
2
44521.8 143
0
9 Terminal~
194 98 647 0 1 3
0 54
0
0 0 49520 90
6 clock0
-48 -4 -6 4
2 T4
-7 -32 7 -24
0
7 clock0;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9513 0 0
2
44521.8 144
0
9 Terminal~
194 98 638 0 1 3
0 53
0
0 0 49520 90
6 clock1
-45 -6 -3 2
2 T3
-7 -32 7 -24
0
7 clock1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4896 0 0
2
44521.8 145
0
9 Terminal~
194 282 559 0 1 3
0 54
0
0 0 49520 270
6 clock0
2 -5 44 3
2 T2
-7 -32 7 -24
0
7 clock0;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4582 0 0
2
44521.8 146
0
9 Terminal~
194 282 550 0 1 3
0 53
0
0 0 49520 270
6 clock1
2 -4 44 4
2 T1
-7 -32 7 -24
0
7 clock1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4121 0 0
2
44521.8 147
0
7 Ground~
168 135 721 0 1 3
0 6
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3664 0 0
2
44521.8 148
0
7 Pulser~
4 74 474 0 10 12
0 126 127 17 48 0 0 10 10 8
8
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3124 0 0
2
44521.8 149
0
14 NO PushButton~
191 477 317 0 2 5
0 33 62
0
0 0 4208 0
0
3 S15
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
4395 0 0
2
44521.8 150
0
14 NO PushButton~
191 396 316 0 2 5
0 34 62
0
0 0 4208 0
0
3 S14
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
4729 0 0
2
44521.8 151
0
14 NO PushButton~
191 314 316 0 2 5
0 35 62
0
0 0 4208 0
0
3 S13
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3472 0 0
2
44521.8 152
0
14 NO PushButton~
191 478 254 0 2 5
0 33 65
0
0 0 4208 0
0
3 S11
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
9236 0 0
2
44521.8 153
0
14 NO PushButton~
191 397 253 0 2 5
0 34 65
0
0 0 4208 0
0
3 S10
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
9829 0 0
2
44521.8 154
0
14 NO PushButton~
191 315 253 0 2 5
0 35 65
0
0 0 4208 0
0
2 S9
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
8397 0 0
2
44521.8 155
0
14 NO PushButton~
191 478 191 0 2 5
0 33 64
0
0 0 4208 0
0
2 S7
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3297 0 0
2
44521.8 156
0
14 NO PushButton~
191 397 190 0 2 5
0 34 64
0
0 0 4208 0
0
2 S5
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
6696 0 0
2
44521.8 157
0
14 NO PushButton~
191 315 190 0 2 5
0 35 64
0
0 0 4208 0
0
2 S4
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
8438 0 0
2
44521.8 158
0
14 NO PushButton~
191 477 128 0 2 5
0 33 63
0
0 0 4208 0
0
2 S3
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3768 0 0
2
44521.8 159
0
14 NO PushButton~
191 396 127 0 2 5
0 34 63
0
0 0 4208 0
0
2 S2
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
9851 0 0
2
44521.8 160
0
14 NO PushButton~
191 314 127 0 2 5
0 35 63
0
0 0 4208 0
0
2 S1
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
5881 0 0
2
44521.8 161
0
9 Resistor~
219 2309 136 0 4 5
0 41 6 0 -1
0
0 0 880 90
2 1k
8 0 22 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9387 0 0
2
44521.8 162
0
9 Resistor~
219 433 90 0 4 5
0 34 93 0 1
0
0 0 880 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3321 0 0
2
44521.8 163
0
9 Resistor~
219 514 89 0 4 5
0 33 93 0 1
0
0 0 880 90
2 1k
8 0 22 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5764 0 0
2
44521.8 164
0
9 Resistor~
219 343 89 0 4 5
0 35 93 0 1
0
0 0 880 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3559 0 0
2
44521.8 165
0
305
1 4 2 0 0 4112 0 3 53 0 0 2
1156 300
1156 261
1 1 3 0 0 0 0 4 5 0 0 2
822 289
822 289
1 1 4 0 0 4096 0 7 6 0 0 2
939 287
939 290
1 1 5 0 0 4224 0 1 8 0 0 2
658 107
696 107
2 1 6 0 0 8192 0 274 9 0 0 4
2309 118
2309 103
2355 103
2355 115
1 0 41 0 0 4096 0 274 0 0 79 3
2309 154
2309 177
2308 177
1 0 8 0 0 4096 0 11 0 0 32 3
1250 1684
1201 1684
1201 1686
20 0 20 0 0 8192 0 208 0 0 112 3
1710 377
1741 377
1741 217
19 2 66 0 0 8320 0 208 13 0 0 4
1710 368
1729 368
1729 288
1667 288
1 1 7 0 0 4096 0 12 13 0 0 2
1594 288
1631 288
1 0 11 0 0 8320 0 16 0 0 143 3
1608 669
1569 669
1569 566
0 1 10 0 0 4224 0 0 15 144 0 3
1561 557
1561 656
1614 656
0 1 9 0 0 4224 0 0 14 145 0 3
1573 548
1573 644
1620 644
1 3 9 0 0 0 0 18 17 0 0 2
1267 286
1267 261
1 2 10 0 0 0 0 19 17 0 0 2
1273 273
1273 261
1 1 11 0 0 0 0 20 17 0 0 2
1279 261
1279 261
1 1 2 0 0 0 0 25 21 0 0 2
1639 1541
1621 1541
4 1 12 0 0 4224 0 25 22 0 0 2
1639 1568
1621 1568
3 1 13 0 0 4224 0 25 23 0 0 2
1639 1559
1621 1559
2 1 14 0 0 4096 0 25 24 0 0 2
1639 1550
1621 1550
4 1 67 0 0 8320 0 29 27 0 0 4
1431 1634
1440 1634
1440 1712
1464 1712
1 3 15 0 0 4096 0 26 27 0 0 3
1536 1722
1510 1722
1510 1721
1 0 16 0 0 4096 0 28 0 0 25 3
1167 1599
1167 1625
1166 1625
1 0 16 0 0 8192 0 136 0 0 25 3
1123 1664
1111 1664
1111 1625
1 3 16 0 0 4224 0 29 138 0 0 2
1386 1625
1106 1625
1 0 6 0 0 12288 0 35 0 0 27 4
935 1237
935 1226
909 1226
909 1309
4 1 6 0 0 0 0 35 30 0 0 4
935 1300
935 1309
900 1309
900 1314
1 3 17 0 0 4096 0 31 35 0 0 2
895 1276
911 1276
2 3 68 0 0 4224 0 35 34 0 0 2
911 1258
868 1258
1 2 18 0 0 4096 0 32 34 0 0 2
793 1267
822 1267
1 1 19 0 0 4096 0 33 34 0 0 2
792 1249
822 1249
2 0 8 0 0 12416 0 27 0 0 100 5
1464 1730
1341 1730
1341 1698
1201 1698
1201 1673
3 2 69 0 0 8320 0 29 37 0 0 3
1386 1643
1376 1643
1376 1659
1 1 4 0 0 12288 0 37 38 0 0 4
1376 1695
1376 1694
1376 1694
1376 1711
1 1 20 0 0 0 0 40 39 0 0 2
1299 1634
1329 1634
2 2 70 0 0 4224 0 39 29 0 0 2
1365 1634
1386 1634
1 1 21 0 0 4096 0 41 42 0 0 2
1091 354
1160 354
0 1 21 0 0 0 0 0 43 207 0 3
2435 186
2435 143
2436 143
1 1 22 0 0 8192 0 44 2 0 0 3
1150 95
1150 96
1114 96
1 3 22 0 0 4224 0 45 113 0 0 3
1586 929
1586 1015
1603 1015
1 3 14 0 0 4224 0 52 53 0 0 2
1162 286
1162 261
1 2 13 0 0 0 0 51 53 0 0 2
1168 273
1168 261
1 1 12 0 0 0 0 50 53 0 0 2
1174 261
1174 261
1 3 23 0 0 4096 0 47 46 0 0 2
1078 288
1078 263
1 2 24 0 0 4096 0 48 46 0 0 2
1084 275
1084 263
1 1 25 0 0 0 0 49 46 0 0 2
1090 263
1090 263
1 3 26 0 0 4096 0 54 55 0 0 2
912 118
912 113
1 4 29 0 0 4096 0 58 55 0 0 2
906 118
906 113
1 2 28 0 0 4096 0 57 55 0 0 2
918 118
918 113
1 1 27 0 0 4096 0 56 55 0 0 2
924 118
924 113
2 1 18 0 0 4096 0 61 59 0 0 2
924 773
973 773
1 1 71 0 0 8320 0 69 60 0 0 3
774 755
758 755
758 733
0 1 30 0 0 8192 0 0 62 55 0 3
862 773
862 732
906 732
1 11 6 0 0 0 0 63 69 0 0 3
852 792
852 755
844 755
13 1 30 0 0 4224 0 69 61 0 0 2
838 773
888 773
1 5 31 0 0 4096 0 64 69 0 0 2
752 791
774 791
1 6 32 0 0 4096 0 65 69 0 0 2
752 800
774 800
1 2 33 0 0 4096 0 66 69 0 0 2
752 764
774 764
1 3 34 0 0 4096 0 67 69 0 0 2
752 773
774 773
1 4 35 0 0 4096 0 68 69 0 0 2
752 782
774 782
0 0 72 0 0 4224 0 0 0 0 0 5
595 393
1013 393
1013 32
595 32
595 393
1 0 19 0 0 0 0 77 0 0 63 2
1669 185
1669 168
1 3 19 0 0 0 0 78 79 0 0 3
1669 153
1669 168
1659 168
2 1 36 0 0 8192 0 79 80 0 0 3
1614 177
1598 177
1598 200
2 1 73 0 0 4224 0 75 79 0 0 2
1604 159
1614 159
1 1 18 0 0 4224 0 76 36 0 0 2
1664 69
1557 69
1 1 5 0 0 0 0 74 75 0 0 2
1554 159
1568 159
1 -208000 37 0 0 4096 0 81 0 0 199 2
2119 465
2062 465
1 -207999 38 0 0 4096 0 82 0 0 199 2
2119 451
2062 451
1 -207998 39 0 0 4096 0 83 0 0 199 2
2119 435
2062 435
1 -207997 40 0 0 4096 0 84 0 0 199 2
2119 417
2062 417
14 1 37 0 0 0 0 241 86 0 0 2
816 614
831 614
13 1 38 0 0 0 0 241 85 0 0 2
816 596
831 596
12 1 39 0 0 0 0 241 87 0 0 2
816 578
831 578
11 1 40 0 0 0 0 241 88 0 0 2
816 560
831 560
0 1 36 0 0 4224 0 0 89 113 0 2
1702 1553
1779 1553
1 3 7 0 0 4096 0 10 92 0 0 2
2285 195
2337 195
1 2 20 0 0 0 0 90 92 0 0 2
2285 186
2337 186
1 1 41 0 0 4096 0 91 92 0 0 2
2284 177
2337 177
2 1 43 0 0 4096 0 202 94 0 0 2
2514 479
2488 479
1 2 42 0 0 4096 0 93 205 0 0 2
2485 619
2517 619
1 2 44 0 0 4096 0 95 199 0 0 2
2484 331
2514 331
-3260 1 41 0 0 4096 0 0 97 226 0 2
1823 481
1879 481
1 -3264 42 0 0 4096 0 99 0 0 226 2
1880 550
1823 550
1 -3262 44 0 0 4096 0 100 0 0 226 2
1880 519
1823 519
1 -3263 43 0 0 4096 0 98 0 0 226 2
1880 535
1823 535
1 -3261 45 0 0 4096 0 101 0 0 226 2
1880 504
1823 504
1 1 6 0 0 12288 0 104 107 0 0 4
1967 1243
1967 1229
1936 1229
1936 1320
2 1 74 0 0 4224 0 104 106 0 0 3
1943 1264
1920 1264
1920 1249
1 4 8 0 0 0 0 105 104 0 0 2
1967 1318
1967 1306
6 1 20 0 0 0 0 104 102 0 0 3
1991 1264
2049 1264
2049 1263
3 1 19 0 0 4224 0 104 103 0 0 3
1943 1282
1901 1282
1901 1281
14 -3260 41 0 0 4224 0 208 0 0 226 2
1704 413
1823 413
4 -3260 41 0 0 0 0 206 0 0 226 2
1927 312
1823 312
12 1 75 0 0 4224 0 206 108 0 0 3
1991 312
2026 312
2026 277
1 1 6 0 0 0 0 176 109 0 0 4
1710 1238
1710 1224
1679 1224
1679 1315
2 1 76 0 0 4224 0 176 110 0 0 3
1686 1259
1663 1259
1663 1244
1 4 46 0 0 4096 0 111 176 0 0 2
1710 1313
1710 1301
1 2 77 0 0 4224 0 112 190 0 0 3
1293 955
1293 1007
1342 1007
1 3 8 0 0 0 0 134 136 0 0 2
1220 1673
1168 1673
1 0 6 0 0 0 0 113 0 0 107 3
1603 997
1592 997
1592 1033
1 2 15 0 0 4224 0 120 113 0 0 2
1578 1006
1609 1006
1 4 20 0 0 0 0 119 113 0 0 2
1578 1024
1609 1024
8 0 6 0 0 0 0 113 0 0 107 2
1609 1060
1592 1060
7 0 6 0 0 0 0 113 0 0 107 2
1609 1051
1592 1051
6 0 6 0 0 0 0 113 0 0 107 2
1609 1042
1592 1042
5 1 6 0 0 0 0 113 118 0 0 3
1609 1033
1592 1033
1592 1111
1 12 14 0 0 0 0 114 113 0 0 2
1687 1042
1673 1042
1 11 2 0 0 4224 0 117 113 0 0 2
1739 1033
1673 1033
1 14 12 0 0 0 0 116 113 0 0 2
1687 1060
1673 1060
1 13 13 0 0 0 0 115 113 0 0 2
1687 1051
1673 1051
1 18 20 0 0 12416 0 121 206 0 0 6
1762 154
1741 154
1741 217
2007 217
2007 276
1991 276
2 5 36 0 0 0 0 127 25 0 0 4
1713 1532
1702 1532
1702 1554
1689 1554
1 3 47 0 0 4096 0 126 127 0 0 2
1796 1523
1758 1523
1 1 48 0 0 4096 0 127 128 0 0 2
1713 1514
1690 1514
1 3 46 0 0 4224 0 125 123 0 0 2
1795 1467
1757 1467
1 2 7 0 0 0 0 124 123 0 0 2
1690 1476
1712 1476
1 1 20 0 0 0 0 123 122 0 0 2
1712 1458
1689 1458
6 3 78 0 0 4224 0 164 132 0 0 3
1491 557
1276 557
1276 604
1 0 79 0 0 4096 0 132 0 0 154 2
1267 649
1267 656
1 1 14 0 0 0 0 130 131 0 0 2
1276 730
1276 711
1 2 2 0 0 0 0 129 131 0 0 2
1294 731
1294 711
2 3 80 0 0 4224 0 132 131 0 0 2
1285 649
1285 665
2 3 81 0 0 4224 0 133 190 0 0 4
1396 962
1311 962
1311 1016
1336 1016
11 1 82 0 0 8320 0 190 133 0 0 4
1406 1034
1446 1034
1446 962
1432 962
1 2 20 0 0 0 0 135 136 0 0 2
1047 1682
1123 1682
1 1 7 0 0 0 0 137 138 0 0 2
1045 1616
1061 1616
1 2 48 0 0 0 0 139 138 0 0 2
1045 1634
1061 1634
14 1 51 0 0 4096 0 146 142 0 0 2
219 690
221 690
13 1 52 0 0 4096 0 146 143 0 0 2
219 681
221 681
12 1 50 0 0 4224 0 146 141 0 0 2
219 672
221 672
11 1 49 0 0 4224 0 146 140 0 0 2
219 663
221 663
6 0 6 0 0 0 0 146 0 0 300 2
143 690
135 690
1 5 54 0 0 4096 0 145 146 0 0 2
107 681
149 681
1 4 53 0 0 4096 0 144 146 0 0 2
107 672
149 672
10 1 63 0 0 4096 0 146 253 0 0 2
219 654
221 654
9 1 64 0 0 4096 0 146 252 0 0 2
219 645
221 645
8 1 65 0 0 4096 0 146 254 0 0 2
219 636
221 636
7 1 62 0 0 4096 0 146 255 0 0 2
219 627
221 627
10 -1535 11 0 0 0 0 208 0 0 146 2
1640 449
1596 449
9 -1534 10 0 0 0 0 208 0 0 146 2
1640 440
1596 440
8 -1533 9 0 0 0 0 208 0 0 146 2
1640 431
1596 431
13 -1535 11 0 0 0 0 164 0 0 146 2
1555 566
1596 566
12 -1534 10 0 0 0 0 164 0 0 146 2
1555 557
1596 557
11 -1533 9 0 0 0 0 164 0 0 146 2
1555 548
1596 548
-95129 0 1 0 0 4128 0 0 0 0 0 2
1596 352
1596 624
0 1 79 0 0 4096 0 0 154 154 0 3
1331 656
1403 656
1403 651
1 2 2 0 0 0 0 157 155 0 0 2
1430 728
1430 712
1 1 12 0 0 0 0 156 155 0 0 2
1412 728
1412 712
2 3 83 0 0 4224 0 154 155 0 0 2
1421 651
1421 666
1 2 2 0 0 0 0 153 149 0 0 2
1358 726
1358 710
1 1 13 0 0 0 0 152 149 0 0 2
1340 726
1340 710
1 1 20 0 0 0 0 148 151 0 0 2
1175 656
1206 656
2 1 79 0 0 4224 0 151 150 0 0 3
1242 656
1331 656
1331 649
2 3 84 0 0 4224 0 150 149 0 0 2
1349 649
1349 664
3 7 85 0 0 8320 0 150 164 0 0 3
1340 604
1340 566
1491 566
7 0 6 0 0 0 0 208 0 0 232 2
1640 422
1624 422
1 14 25 0 0 4096 0 160 190 0 0 2
1419 1061
1406 1061
1 13 24 0 0 4096 0 159 190 0 0 2
1419 1052
1406 1052
1 12 23 0 0 0 0 158 190 0 0 2
1419 1043
1406 1043
14 0 6 0 0 0 0 164 0 0 168 4
1555 593
1565 593
1565 611
1475 611
1 2 23 0 0 4224 0 161 164 0 0 2
1458 521
1491 521
1 3 24 0 0 4224 0 162 164 0 0 2
1458 530
1491 530
1 4 25 0 0 4224 0 163 164 0 0 2
1458 539
1491 539
3 8 86 0 0 8320 0 154 164 0 0 3
1412 606
1412 575
1491 575
9 0 6 0 0 0 0 164 0 0 168 2
1491 593
1475 593
5 0 6 0 0 0 0 164 0 0 168 2
1491 548
1475 548
1 1 6 0 0 8320 0 164 165 0 0 3
1491 512
1475 512
1475 658
4 1 48 0 0 4096 0 261 168 0 0 4
104 474
129 474
129 485
154 485
2 2 87 0 0 4224 0 169 167 0 0 2
1347 1504
1363 1504
3 1 55 0 0 4096 0 167 170 0 0 2
1408 1495
1452 1495
1 1 2 0 0 0 0 171 169 0 0 3
1267 1502
1267 1504
1311 1504
1 1 48 0 0 4224 0 167 172 0 0 2
1363 1486
1304 1486
3 1 56 0 0 4096 0 166 175 0 0 2
1103 1495
1134 1495
1 2 2 0 0 0 0 174 166 0 0 3
1035 1503
1035 1504
1058 1504
1 1 17 0 0 4224 0 166 173 0 0 2
1058 1486
1000 1486
6 1 3 0 0 4224 0 176 178 0 0 3
1734 1259
1792 1259
1792 1258
3 1 47 0 0 4224 0 176 177 0 0 3
1686 1277
1644 1277
1644 1276
1 1 6 0 0 0 0 179 184 0 0 4
1400 1238
1400 1220
1371 1220
1371 1331
6 1 4 0 0 4224 0 179 183 0 0 3
1424 1259
1482 1259
1482 1258
1 4 55 0 0 4224 0 182 179 0 0 3
1332 1313
1400 1313
1400 1301
3 1 56 0 0 4224 0 179 181 0 0 3
1376 1277
1299 1277
1299 1275
1 2 88 0 0 8320 0 180 179 0 0 3
1339 1256
1339 1259
1376 1259
1 1 6 0 0 0 0 189 185 0 0 4
1105 1239
1105 1221
1076 1221
1076 1332
6 1 7 0 0 4224 0 189 186 0 0 3
1129 1260
1187 1260
1187 1259
1 4 16 0 0 0 0 187 189 0 0 3
1037 1314
1105 1314
1105 1302
3 6 89 0 0 4224 0 189 35 0 0 4
1081 1278
985 1278
985 1258
959 1258
1 2 90 0 0 8320 0 188 189 0 0 3
1044 1257
1044 1260
1081 1260
1 1 8 0 0 0 0 190 192 0 0 2
1342 998
1260 998
0 4 6 0 0 0 0 0 190 194 0 3
1326 1034
1326 1025
1342 1025
8 0 6 0 0 0 0 190 0 0 194 2
1342 1061
1325 1061
7 0 6 0 0 0 0 190 0 0 194 2
1342 1052
1325 1052
6 0 6 0 0 0 0 190 0 0 194 2
1342 1043
1325 1043
5 1 6 0 0 0 0 190 191 0 0 3
1342 1034
1325 1034
1325 1107
13 -207997 40 0 0 4224 0 206 0 0 199 2
1991 321
2062 321
14 -207998 39 0 0 4224 0 206 0 0 199 2
1991 330
2062 330
15 -207999 38 0 0 4224 0 206 0 0 199 2
1991 339
2062 339
16 -208000 37 0 0 4224 0 206 0 0 199 2
1991 348
2062 348
-13308169 0 1 0 0 4256 0 0 0 0 0 2
2062 138
2062 707
1 17 6 0 0 0 0 193 206 0 0 3
1904 296
1904 276
1921 276
5 -3261 45 0 0 4096 0 206 0 0 226 2
1927 321
1823 321
6 -3262 44 0 0 4096 0 206 0 0 226 2
1927 330
1823 330
7 -3263 43 0 0 4096 0 206 0 0 226 2
1927 339
1823 339
3 0 21 0 0 4096 0 194 0 0 207 2
2517 207
2435 207
3 0 21 0 0 0 0 199 0 0 207 2
2514 349
2435 349
3 0 21 0 0 0 0 202 0 0 207 2
2514 497
2435 497
4 3 21 0 0 8320 0 92 205 0 0 4
2382 186
2435 186
2435 637
2517 637
6 1 27 0 0 4224 0 205 70 0 0 2
2565 619
2612 619
4 1 6 0 0 0 0 205 203 0 0 2
2541 661
2541 673
1 1 6 0 0 0 0 205 204 0 0 4
2541 598
2541 559
2641 559
2641 572
6 1 28 0 0 4224 0 202 71 0 0 2
2562 479
2608 479
4 1 6 0 0 0 0 202 200 0 0 2
2538 521
2538 533
1 1 6 0 0 0 0 202 201 0 0 4
2538 458
2538 419
2645 419
2645 428
6 1 26 0 0 4224 0 199 72 0 0 3
2562 331
2611 331
2611 332
4 1 6 0 0 0 0 199 197 0 0 2
2538 373
2538 387
1 1 6 0 0 0 0 199 198 0 0 4
2538 310
2538 273
2645 273
2645 284
6 1 29 0 0 4224 0 194 73 0 0 2
2565 189
2613 189
4 1 6 0 0 0 0 194 196 0 0 2
2541 231
2541 243
1 1 6 0 0 0 0 194 195 0 0 4
2541 168
2541 129
2647 129
2647 143
1 2 45 0 0 0 0 96 194 0 0 2
2487 189
2517 189
8 -3264 42 0 0 4096 0 206 0 0 226 2
1927 348
1823 348
15 -3261 45 0 0 4224 0 208 0 0 226 2
1704 422
1823 422
16 -3262 44 0 0 4224 0 208 0 0 226 2
1704 431
1823 431
17 -3263 43 0 0 4224 0 208 0 0 226 2
1704 440
1823 440
18 -3264 42 0 0 4224 0 208 0 0 226 2
1704 449
1823 449
-846037834 0 1 0 0 32 0 0 0 0 0 2
1823 140
1823 709
6 0 6 0 0 0 0 208 0 0 232 2
1640 413
1624 413
5 0 6 0 0 0 0 208 0 0 232 2
1640 404
1624 404
4 0 6 0 0 0 0 208 0 0 232 2
1640 395
1624 395
3 0 6 0 0 0 0 208 0 0 232 2
1640 386
1624 386
2 0 6 0 0 0 0 208 0 0 232 2
1640 377
1624 377
1 1 6 0 0 0 0 208 207 0 0 3
1640 368
1624 368
1624 473
0 1 61 0 0 8192 0 0 226 250 0 3
555 721
555 730
572 730
2 0 6 0 0 0 0 209 0 0 241 2
515 542
506 542
4 1 32 0 0 0 0 209 215 0 0 2
515 560
494 560
1 3 31 0 0 0 0 220 209 0 0 2
494 551
515 551
1 13 59 0 0 4224 0 218 209 0 0 2
604 587
579 587
1 12 60 0 0 4224 0 219 209 0 0 2
604 578
579 578
1 11 58 0 0 4224 0 217 209 0 0 2
604 569
579 569
1 10 57 0 0 4224 0 216 209 0 0 2
604 560
579 560
1 0 6 0 0 0 0 209 0 0 243 3
515 533
506 533
506 569
9 0 6 0 0 0 0 209 0 0 243 2
515 614
506 614
5 1 6 0 0 0 0 209 214 0 0 3
515 569
506 569
506 629
1 8 52 0 0 4224 0 213 209 0 0 2
500 596
515 596
2 7 91 0 0 4224 0 210 209 0 0 2
441 587
515 587
1 1 50 0 0 0 0 212 210 0 0 2
404 587
405 587
1 6 51 0 0 4224 0 211 209 0 0 2
500 578
515 578
1 1 32 0 0 0 0 221 222 0 0 2
494 721
501 721
1 1 31 0 0 4096 0 225 227 0 0 2
572 739
546 739
1 2 61 0 0 4224 0 224 222 0 0 2
572 721
537 721
1 0 61 0 0 0 0 223 0 0 250 3
572 712
548 712
548 721
0 1 17 0 0 0 0 0 228 254 0 2
117 465
154 465
3 3 92 0 0 4224 0 229 147 0 0 2
126 549
153 549
1 3 17 0 0 0 0 229 261 0 0 6
81 540
63 540
63 514
117 514
117 465
98 465
1 2 30 0 0 0 0 230 229 0 0 2
69 558
81 558
1 1 62 0 0 0 0 231 241 0 0 2
752 542
752 542
1 8 59 0 0 0 0 233 241 0 0 2
752 605
752 605
1 9 31 0 0 0 0 232 241 0 0 2
752 614
752 614
1 6 60 0 0 0 0 235 241 0 0 4
752 587
753 587
753 587
752 587
1 7 61 0 0 0 0 234 241 0 0 2
752 596
752 596
1 4 58 0 0 0 0 237 241 0 0 2
752 569
752 569
1 5 61 0 0 0 0 236 241 0 0 2
752 578
752 578
1 2 57 0 0 0 0 239 241 0 0 2
752 551
752 551
1 3 61 0 0 0 0 238 241 0 0 2
752 560
752 560
1 10 6 0 0 0 0 240 241 0 0 3
739 639
739 623
746 623
6 1 32 0 0 4224 0 147 246 0 0 2
223 540
270 540
5 1 31 0 0 4224 0 147 245 0 0 2
223 531
270 531
2 0 6 0 0 0 0 147 0 0 269 2
159 540
135 540
0 1 6 0 0 0 0 0 147 300 0 3
135 654
135 531
159 531
2 0 63 0 0 4096 0 273 0 0 299 2
297 135
297 153
2 0 63 0 0 0 0 272 0 0 299 2
379 135
379 153
2 0 64 0 0 4096 0 270 0 0 298 2
298 198
298 216
2 0 64 0 0 0 0 269 0 0 298 2
380 198
380 216
2 0 65 0 0 4096 0 267 0 0 297 2
298 261
298 279
2 0 65 0 0 0 0 266 0 0 297 2
380 261
380 279
2 0 62 0 0 4096 0 264 0 0 296 2
297 324
297 342
2 0 62 0 0 0 0 263 0 0 296 2
379 324
379 342
1 0 33 0 0 0 0 262 0 0 292 2
494 325
514 325
1 0 33 0 0 0 0 265 0 0 292 2
495 262
514 262
1 0 33 0 0 0 0 268 0 0 292 2
495 199
514 199
1 0 34 0 0 0 0 263 0 0 293 2
413 324
433 324
1 0 34 0 0 0 0 266 0 0 293 2
414 261
433 261
1 0 34 0 0 0 0 269 0 0 293 2
414 198
433 198
1 0 35 0 0 0 0 264 0 0 294 2
331 324
343 324
1 0 35 0 0 0 0 267 0 0 294 2
332 261
343 261
1 0 35 0 0 0 0 270 0 0 294 2
332 198
343 198
1 0 33 0 0 0 0 271 0 0 292 2
494 136
514 136
1 0 34 0 0 0 0 272 0 0 293 2
413 135
433 135
1 0 35 0 0 0 0 273 0 0 294 2
331 135
343 135
2 2 93 0 0 8192 0 275 276 0 0 3
433 72
433 71
514 71
2 2 93 0 0 4224 0 277 275 0 0 3
343 71
433 71
433 72
1 1 33 0 0 4224 0 276 242 0 0 2
514 107
514 351
1 1 34 0 0 4224 0 275 243 0 0 2
433 108
433 353
1 1 35 0 0 4224 0 277 244 0 0 2
343 107
343 388
2 1 93 0 0 0 0 277 247 0 0 2
343 71
343 64
1 2 62 0 0 4224 0 251 262 0 0 3
216 342
460 342
460 325
1 2 65 0 0 4224 0 250 265 0 0 3
215 279
461 279
461 262
1 2 64 0 0 4224 0 249 268 0 0 3
217 216
461 216
461 199
1 2 63 0 0 4224 0 248 271 0 0 3
217 153
460 153
460 136
3 1 6 0 0 0 0 146 260 0 0 3
143 654
135 654
135 715
1 2 54 0 0 0 0 256 146 0 0 2
109 645
149 645
1 1 53 0 0 0 0 257 146 0 0 2
109 636
149 636
0 1 54 0 0 0 0 0 258 305 0 2
234 558
270 558
7 1 53 0 0 4224 0 147 259 0 0 2
223 549
270 549
8 4 54 0 0 12416 0 147 147 0 0 6
223 558
234 558
234 575
144 575
144 558
153 558
43
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 26
616 156 719 220
623 161 711 209
26      INPUTS

<-- teclado
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
780 312 883 336
787 317 875 333
11 DDispon�vel
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
920 313 991 337
927 319 983 335
7 Overrun
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
887 157 942 181
894 162 934 178
5 SAIDA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 222
905 1745 1314 1892
913 1752 1305 1872
222 IF !clock AND write_read_out:
   write_read = 0
   IF (modo==0 AND overrun=0):  // escrita
      q += 1
   ELSE:          // leitura
      q -= 1      // (feito pelo pq acima tamb�m)
      inicio += 1
      modo = 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
1227 172 1306 196
1234 177 1298 193
8 endereco
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
2031 1313 2074 1357
2036 1317 2068 1349
4 modo
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
1720 1325 1823 1349
1727 1330 1815 1346
11 ddisponivel
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1401 1323 1472 1347
1408 1329 1464 1345
7 overrun
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1342 1080 1405 1104
1349 1086 1397 1102
6 inicio
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
64 73 119 97
71 78 111 94
5 saida
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 24
437 672 640 696
442 676 634 692
24 aritmetica para *, 0 e #
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
454 479 617 503
459 483 611 499
19 aritmetica para 1-9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
147 428 282 452
150 430 278 446
16 divisao do clock
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
299 288 330 312
302 290 326 306
3 (*)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
462 289 493 313
465 291 489 307
3 (#)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
381 288 412 312
384 290 408 306
3 (0)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
463 226 494 250
466 228 490 244
3 (9)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
382 225 413 249
385 227 409 243
3 (8)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
300 225 331 249
303 227 327 243
3 (7)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
463 163 494 187
466 165 490 181
3 (6)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
382 162 413 186
385 164 409 180
3 (5)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
300 162 331 186
303 164 327 180
3 (4)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
462 99 493 123
465 101 489 117
3 (3)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
381 98 412 122
384 100 408 116
3 (2)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
295 93 334 117
302 99 326 115
3 (1)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
397 37 540 61
404 42 532 58
16 matriz de botoes
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
55 93 120 132
63 100 111 130
14 * -> E
# -> F
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
958 1326 1053 1350
965 1331 1045 1347
10 write/read
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 24
1016 1521 1139 1565
1021 1525 1133 1557
24 clock AND q=8:
   or_up
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 32
1292 1522 1463 1566
1297 1526 1457 1558
32 clock_down AND q!=8:
   or_down
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 103
1254 411 1465 535
1259 415 1459 511
103 ESCRITA (modo=0)
end = inicio + 7 (se q=8)
    = inicio + q (senao)

LEITURA (modo=1)
end = inicio
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
1601 1087 1696 1111
1608 1092 1688 1108
10 quantidade
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 154
1856 1459 2423 1563
1863 1465 2415 1545
154 IF write_read AND (modo == 1):  // operacao no clockup
   ddown = 1

IF nclock AND (q > 0):  // operacao no clockup (pr�ximo ap�s mudar q)
   ddup = 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1428 52 1491 76
1435 57 1483 73
6 insert
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1431 138 1478 162
1438 144 1470 160
4 read
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
2711 338 2814 362
2718 343 2806 359
11 REGISTRADOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 51
675 450 842 514
682 455 834 503
51 multiplex para
escolher entre
as duas aritmeticas
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
749 866 916 890
756 871 908 887
19 controle das teclas
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
611 55 682 79
618 60 674 76
7 leTecla
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
1122 172 1217 196
1129 177 1209 193
10 quantidade
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1048 172 1111 196
1055 178 1103 194
6 inicio
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
1107 140 1202 164
1114 145 1194 161
10 para debug
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-06 1e-07 1e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
